
module LCD_CTRL_DW01_add_5 ( A, B, CI, SUM, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [9:1] carry;

  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(SUM[8]), .S(SUM[7]) );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module LCD_CTRL_DW01_add_4 ( A, B, CI, SUM, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [9:1] carry;

  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFHX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  CMPR32X2 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(A[8]), .B(carry[8]), .Y(SUM[8]) );
  AND2X2 U3 ( .A(A[8]), .B(carry[8]), .Y(SUM[9]) );
  XOR2X1 U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module LCD_CTRL_DW01_add_3 ( A, B, CI, SUM, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6;
  wire   [9:1] carry;

  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFHX4 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFHX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  XOR2X4 U1 ( .A(B[9]), .B(n5), .Y(SUM[9]) );
  XOR2XL U2 ( .A(B[5]), .B(A[5]), .Y(n1) );
  XOR2XL U3 ( .A(carry[5]), .B(n1), .Y(SUM[5]) );
  NAND2X1 U4 ( .A(B[5]), .B(carry[5]), .Y(n2) );
  NAND2X1 U5 ( .A(A[5]), .B(carry[5]), .Y(n3) );
  NAND2XL U6 ( .A(A[5]), .B(B[5]), .Y(n4) );
  NAND3X1 U7 ( .A(n2), .B(n3), .C(n4), .Y(carry[6]) );
  XOR2X1 U8 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  AND2X2 U9 ( .A(B[8]), .B(carry[8]), .Y(n5) );
  OAI2BB1X1 U10 ( .A0N(A[1]), .A1N(B[1]), .B0(n6), .Y(carry[2]) );
  OAI211X1 U11 ( .A0(A[1]), .A1(B[1]), .B0(A[0]), .C0(B[0]), .Y(n6) );
endmodule


module LCD_CTRL ( clk, reset, cmd, cmd_valid, IROM_Q, IROM_rd, IROM_A, 
        IRAM_valid, IRAM_D, IRAM_A, busy, done );
  input [3:0] cmd;
  input [7:0] IROM_Q;
  output [5:0] IROM_A;
  output [7:0] IRAM_D;
  output [5:0] IRAM_A;
  input clk, reset, cmd_valid;
  output IROM_rd, IRAM_valid, busy, done;
  wire   N2484, N2485, N2486, N2488, N2489, N2490, N2491, N2492, N2493, N2494,
         N2495, N2497, N2498, N2501, N2502, N2503, N2504, N2505, N2506, N2507,
         N2508, N2509, N2510, N2512, N2513, N2514, N2515, N2516, N2517, N2518,
         N2519, N2520, N2521, N2522, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, \state_cs[0] ,
         N2538, N2541, N2545, N2546, N2547, N2548, N2549, N2568, N2569, N2570,
         N2571, N2572, N2613, N2614, N2615, N2617, N2623, N2624, N2625, N2630,
         N2631, N2632, N2633, N2634, N2635, \ImageBuffer[63][7] ,
         \ImageBuffer[63][6] , \ImageBuffer[63][5] , \ImageBuffer[63][4] ,
         \ImageBuffer[63][3] , \ImageBuffer[63][2] , \ImageBuffer[63][1] ,
         \ImageBuffer[63][0] , \ImageBuffer[62][7] , \ImageBuffer[62][6] ,
         \ImageBuffer[62][5] , \ImageBuffer[62][4] , \ImageBuffer[62][3] ,
         \ImageBuffer[62][2] , \ImageBuffer[62][1] , \ImageBuffer[62][0] ,
         \ImageBuffer[61][7] , \ImageBuffer[61][6] , \ImageBuffer[61][5] ,
         \ImageBuffer[61][4] , \ImageBuffer[61][3] , \ImageBuffer[61][2] ,
         \ImageBuffer[61][1] , \ImageBuffer[61][0] , \ImageBuffer[60][7] ,
         \ImageBuffer[60][6] , \ImageBuffer[60][5] , \ImageBuffer[60][4] ,
         \ImageBuffer[60][3] , \ImageBuffer[60][2] , \ImageBuffer[60][1] ,
         \ImageBuffer[60][0] , \ImageBuffer[59][7] , \ImageBuffer[59][6] ,
         \ImageBuffer[59][5] , \ImageBuffer[59][4] , \ImageBuffer[59][3] ,
         \ImageBuffer[59][2] , \ImageBuffer[59][1] , \ImageBuffer[59][0] ,
         \ImageBuffer[58][7] , \ImageBuffer[58][6] , \ImageBuffer[58][5] ,
         \ImageBuffer[58][4] , \ImageBuffer[58][3] , \ImageBuffer[58][2] ,
         \ImageBuffer[58][1] , \ImageBuffer[58][0] , \ImageBuffer[57][7] ,
         \ImageBuffer[57][6] , \ImageBuffer[57][5] , \ImageBuffer[57][4] ,
         \ImageBuffer[57][3] , \ImageBuffer[57][2] , \ImageBuffer[57][1] ,
         \ImageBuffer[57][0] , \ImageBuffer[56][7] , \ImageBuffer[56][6] ,
         \ImageBuffer[56][5] , \ImageBuffer[56][4] , \ImageBuffer[56][3] ,
         \ImageBuffer[56][2] , \ImageBuffer[56][1] , \ImageBuffer[56][0] ,
         \ImageBuffer[55][7] , \ImageBuffer[55][6] , \ImageBuffer[55][5] ,
         \ImageBuffer[55][4] , \ImageBuffer[55][3] , \ImageBuffer[55][2] ,
         \ImageBuffer[55][1] , \ImageBuffer[55][0] , \ImageBuffer[54][7] ,
         \ImageBuffer[54][6] , \ImageBuffer[54][5] , \ImageBuffer[54][4] ,
         \ImageBuffer[54][3] , \ImageBuffer[54][2] , \ImageBuffer[54][1] ,
         \ImageBuffer[54][0] , \ImageBuffer[53][7] , \ImageBuffer[53][6] ,
         \ImageBuffer[53][5] , \ImageBuffer[53][4] , \ImageBuffer[53][3] ,
         \ImageBuffer[53][2] , \ImageBuffer[53][1] , \ImageBuffer[53][0] ,
         \ImageBuffer[52][7] , \ImageBuffer[52][6] , \ImageBuffer[52][5] ,
         \ImageBuffer[52][4] , \ImageBuffer[52][3] , \ImageBuffer[52][2] ,
         \ImageBuffer[52][1] , \ImageBuffer[52][0] , \ImageBuffer[51][7] ,
         \ImageBuffer[51][6] , \ImageBuffer[51][5] , \ImageBuffer[51][4] ,
         \ImageBuffer[51][3] , \ImageBuffer[51][2] , \ImageBuffer[51][1] ,
         \ImageBuffer[51][0] , \ImageBuffer[50][7] , \ImageBuffer[50][6] ,
         \ImageBuffer[50][5] , \ImageBuffer[50][4] , \ImageBuffer[50][3] ,
         \ImageBuffer[50][2] , \ImageBuffer[50][1] , \ImageBuffer[50][0] ,
         \ImageBuffer[49][7] , \ImageBuffer[49][6] , \ImageBuffer[49][5] ,
         \ImageBuffer[49][4] , \ImageBuffer[49][3] , \ImageBuffer[49][2] ,
         \ImageBuffer[49][1] , \ImageBuffer[49][0] , \ImageBuffer[48][7] ,
         \ImageBuffer[48][6] , \ImageBuffer[48][5] , \ImageBuffer[48][4] ,
         \ImageBuffer[48][3] , \ImageBuffer[48][2] , \ImageBuffer[48][1] ,
         \ImageBuffer[48][0] , \ImageBuffer[47][7] , \ImageBuffer[47][6] ,
         \ImageBuffer[47][5] , \ImageBuffer[47][4] , \ImageBuffer[47][3] ,
         \ImageBuffer[47][2] , \ImageBuffer[47][1] , \ImageBuffer[47][0] ,
         \ImageBuffer[46][7] , \ImageBuffer[46][6] , \ImageBuffer[46][5] ,
         \ImageBuffer[46][4] , \ImageBuffer[46][3] , \ImageBuffer[46][2] ,
         \ImageBuffer[46][1] , \ImageBuffer[46][0] , \ImageBuffer[45][7] ,
         \ImageBuffer[45][6] , \ImageBuffer[45][5] , \ImageBuffer[45][4] ,
         \ImageBuffer[45][3] , \ImageBuffer[45][2] , \ImageBuffer[45][1] ,
         \ImageBuffer[45][0] , \ImageBuffer[44][7] , \ImageBuffer[44][6] ,
         \ImageBuffer[44][5] , \ImageBuffer[44][4] , \ImageBuffer[44][3] ,
         \ImageBuffer[44][2] , \ImageBuffer[44][1] , \ImageBuffer[44][0] ,
         \ImageBuffer[43][7] , \ImageBuffer[43][6] , \ImageBuffer[43][5] ,
         \ImageBuffer[43][4] , \ImageBuffer[43][3] , \ImageBuffer[43][2] ,
         \ImageBuffer[43][1] , \ImageBuffer[43][0] , \ImageBuffer[42][7] ,
         \ImageBuffer[42][6] , \ImageBuffer[42][5] , \ImageBuffer[42][4] ,
         \ImageBuffer[42][3] , \ImageBuffer[42][2] , \ImageBuffer[42][1] ,
         \ImageBuffer[42][0] , \ImageBuffer[41][7] , \ImageBuffer[41][6] ,
         \ImageBuffer[41][5] , \ImageBuffer[41][4] , \ImageBuffer[41][3] ,
         \ImageBuffer[41][2] , \ImageBuffer[41][1] , \ImageBuffer[41][0] ,
         \ImageBuffer[40][7] , \ImageBuffer[40][6] , \ImageBuffer[40][5] ,
         \ImageBuffer[40][4] , \ImageBuffer[40][3] , \ImageBuffer[40][2] ,
         \ImageBuffer[40][1] , \ImageBuffer[40][0] , \ImageBuffer[39][7] ,
         \ImageBuffer[39][6] , \ImageBuffer[39][5] , \ImageBuffer[39][4] ,
         \ImageBuffer[39][3] , \ImageBuffer[39][2] , \ImageBuffer[39][1] ,
         \ImageBuffer[39][0] , \ImageBuffer[38][7] , \ImageBuffer[38][6] ,
         \ImageBuffer[38][5] , \ImageBuffer[38][4] , \ImageBuffer[38][3] ,
         \ImageBuffer[38][2] , \ImageBuffer[38][1] , \ImageBuffer[38][0] ,
         \ImageBuffer[37][7] , \ImageBuffer[37][6] , \ImageBuffer[37][5] ,
         \ImageBuffer[37][4] , \ImageBuffer[37][3] , \ImageBuffer[37][2] ,
         \ImageBuffer[37][1] , \ImageBuffer[37][0] , \ImageBuffer[36][7] ,
         \ImageBuffer[36][6] , \ImageBuffer[36][5] , \ImageBuffer[36][4] ,
         \ImageBuffer[36][3] , \ImageBuffer[36][2] , \ImageBuffer[36][1] ,
         \ImageBuffer[36][0] , \ImageBuffer[35][7] , \ImageBuffer[35][6] ,
         \ImageBuffer[35][5] , \ImageBuffer[35][4] , \ImageBuffer[35][3] ,
         \ImageBuffer[35][2] , \ImageBuffer[35][1] , \ImageBuffer[35][0] ,
         \ImageBuffer[34][7] , \ImageBuffer[34][6] , \ImageBuffer[34][5] ,
         \ImageBuffer[34][4] , \ImageBuffer[34][3] , \ImageBuffer[34][2] ,
         \ImageBuffer[34][1] , \ImageBuffer[34][0] , \ImageBuffer[33][7] ,
         \ImageBuffer[33][6] , \ImageBuffer[33][5] , \ImageBuffer[33][4] ,
         \ImageBuffer[33][3] , \ImageBuffer[33][2] , \ImageBuffer[33][1] ,
         \ImageBuffer[33][0] , \ImageBuffer[32][7] , \ImageBuffer[32][6] ,
         \ImageBuffer[32][5] , \ImageBuffer[32][4] , \ImageBuffer[32][3] ,
         \ImageBuffer[32][2] , \ImageBuffer[32][1] , \ImageBuffer[32][0] ,
         \ImageBuffer[31][7] , \ImageBuffer[31][6] , \ImageBuffer[31][5] ,
         \ImageBuffer[31][4] , \ImageBuffer[31][3] , \ImageBuffer[31][2] ,
         \ImageBuffer[31][1] , \ImageBuffer[31][0] , \ImageBuffer[30][7] ,
         \ImageBuffer[30][6] , \ImageBuffer[30][5] , \ImageBuffer[30][4] ,
         \ImageBuffer[30][3] , \ImageBuffer[30][2] , \ImageBuffer[30][1] ,
         \ImageBuffer[30][0] , \ImageBuffer[29][7] , \ImageBuffer[29][6] ,
         \ImageBuffer[29][5] , \ImageBuffer[29][4] , \ImageBuffer[29][3] ,
         \ImageBuffer[29][2] , \ImageBuffer[29][1] , \ImageBuffer[29][0] ,
         \ImageBuffer[28][7] , \ImageBuffer[28][6] , \ImageBuffer[28][5] ,
         \ImageBuffer[28][4] , \ImageBuffer[28][3] , \ImageBuffer[28][2] ,
         \ImageBuffer[28][1] , \ImageBuffer[28][0] , \ImageBuffer[27][7] ,
         \ImageBuffer[27][6] , \ImageBuffer[27][5] , \ImageBuffer[27][4] ,
         \ImageBuffer[27][3] , \ImageBuffer[27][2] , \ImageBuffer[27][1] ,
         \ImageBuffer[27][0] , \ImageBuffer[26][7] , \ImageBuffer[26][6] ,
         \ImageBuffer[26][5] , \ImageBuffer[26][4] , \ImageBuffer[26][3] ,
         \ImageBuffer[26][2] , \ImageBuffer[26][1] , \ImageBuffer[26][0] ,
         \ImageBuffer[25][7] , \ImageBuffer[25][6] , \ImageBuffer[25][5] ,
         \ImageBuffer[25][4] , \ImageBuffer[25][3] , \ImageBuffer[25][2] ,
         \ImageBuffer[25][1] , \ImageBuffer[25][0] , \ImageBuffer[24][7] ,
         \ImageBuffer[24][6] , \ImageBuffer[24][5] , \ImageBuffer[24][4] ,
         \ImageBuffer[24][3] , \ImageBuffer[24][2] , \ImageBuffer[24][1] ,
         \ImageBuffer[24][0] , \ImageBuffer[23][7] , \ImageBuffer[23][6] ,
         \ImageBuffer[23][5] , \ImageBuffer[23][4] , \ImageBuffer[23][3] ,
         \ImageBuffer[23][2] , \ImageBuffer[23][1] , \ImageBuffer[23][0] ,
         \ImageBuffer[22][7] , \ImageBuffer[22][6] , \ImageBuffer[22][5] ,
         \ImageBuffer[22][4] , \ImageBuffer[22][3] , \ImageBuffer[22][2] ,
         \ImageBuffer[22][1] , \ImageBuffer[22][0] , \ImageBuffer[21][7] ,
         \ImageBuffer[21][6] , \ImageBuffer[21][5] , \ImageBuffer[21][4] ,
         \ImageBuffer[21][3] , \ImageBuffer[21][2] , \ImageBuffer[21][1] ,
         \ImageBuffer[21][0] , \ImageBuffer[20][7] , \ImageBuffer[20][6] ,
         \ImageBuffer[20][5] , \ImageBuffer[20][4] , \ImageBuffer[20][3] ,
         \ImageBuffer[20][2] , \ImageBuffer[20][1] , \ImageBuffer[20][0] ,
         \ImageBuffer[19][7] , \ImageBuffer[19][6] , \ImageBuffer[19][5] ,
         \ImageBuffer[19][4] , \ImageBuffer[19][3] , \ImageBuffer[19][2] ,
         \ImageBuffer[19][1] , \ImageBuffer[19][0] , \ImageBuffer[18][7] ,
         \ImageBuffer[18][6] , \ImageBuffer[18][5] , \ImageBuffer[18][4] ,
         \ImageBuffer[18][3] , \ImageBuffer[18][2] , \ImageBuffer[18][1] ,
         \ImageBuffer[18][0] , \ImageBuffer[17][7] , \ImageBuffer[17][6] ,
         \ImageBuffer[17][5] , \ImageBuffer[17][4] , \ImageBuffer[17][3] ,
         \ImageBuffer[17][2] , \ImageBuffer[17][1] , \ImageBuffer[17][0] ,
         \ImageBuffer[16][7] , \ImageBuffer[16][6] , \ImageBuffer[16][5] ,
         \ImageBuffer[16][4] , \ImageBuffer[16][3] , \ImageBuffer[16][2] ,
         \ImageBuffer[16][1] , \ImageBuffer[16][0] , \ImageBuffer[15][7] ,
         \ImageBuffer[15][6] , \ImageBuffer[15][5] , \ImageBuffer[15][4] ,
         \ImageBuffer[15][3] , \ImageBuffer[15][2] , \ImageBuffer[15][1] ,
         \ImageBuffer[15][0] , \ImageBuffer[14][7] , \ImageBuffer[14][6] ,
         \ImageBuffer[14][5] , \ImageBuffer[14][4] , \ImageBuffer[14][3] ,
         \ImageBuffer[14][2] , \ImageBuffer[14][1] , \ImageBuffer[14][0] ,
         \ImageBuffer[13][7] , \ImageBuffer[13][6] , \ImageBuffer[13][5] ,
         \ImageBuffer[13][4] , \ImageBuffer[13][3] , \ImageBuffer[13][2] ,
         \ImageBuffer[13][1] , \ImageBuffer[13][0] , \ImageBuffer[12][7] ,
         \ImageBuffer[12][6] , \ImageBuffer[12][5] , \ImageBuffer[12][4] ,
         \ImageBuffer[12][3] , \ImageBuffer[12][2] , \ImageBuffer[12][1] ,
         \ImageBuffer[12][0] , \ImageBuffer[11][7] , \ImageBuffer[11][6] ,
         \ImageBuffer[11][5] , \ImageBuffer[11][4] , \ImageBuffer[11][3] ,
         \ImageBuffer[11][2] , \ImageBuffer[11][1] , \ImageBuffer[11][0] ,
         \ImageBuffer[10][7] , \ImageBuffer[10][6] , \ImageBuffer[10][5] ,
         \ImageBuffer[10][4] , \ImageBuffer[10][3] , \ImageBuffer[10][2] ,
         \ImageBuffer[10][1] , \ImageBuffer[10][0] , \ImageBuffer[9][7] ,
         \ImageBuffer[9][6] , \ImageBuffer[9][5] , \ImageBuffer[9][4] ,
         \ImageBuffer[9][3] , \ImageBuffer[9][2] , \ImageBuffer[9][1] ,
         \ImageBuffer[9][0] , \ImageBuffer[8][7] , \ImageBuffer[8][6] ,
         \ImageBuffer[8][5] , \ImageBuffer[8][4] , \ImageBuffer[8][3] ,
         \ImageBuffer[8][2] , \ImageBuffer[8][1] , \ImageBuffer[8][0] ,
         \ImageBuffer[7][7] , \ImageBuffer[7][6] , \ImageBuffer[7][5] ,
         \ImageBuffer[7][4] , \ImageBuffer[7][3] , \ImageBuffer[7][2] ,
         \ImageBuffer[7][1] , \ImageBuffer[7][0] , \ImageBuffer[6][7] ,
         \ImageBuffer[6][6] , \ImageBuffer[6][5] , \ImageBuffer[6][4] ,
         \ImageBuffer[6][3] , \ImageBuffer[6][2] , \ImageBuffer[6][1] ,
         \ImageBuffer[6][0] , \ImageBuffer[5][7] , \ImageBuffer[5][6] ,
         \ImageBuffer[5][5] , \ImageBuffer[5][4] , \ImageBuffer[5][3] ,
         \ImageBuffer[5][2] , \ImageBuffer[5][1] , \ImageBuffer[5][0] ,
         \ImageBuffer[4][7] , \ImageBuffer[4][6] , \ImageBuffer[4][5] ,
         \ImageBuffer[4][4] , \ImageBuffer[4][3] , \ImageBuffer[4][2] ,
         \ImageBuffer[4][1] , \ImageBuffer[4][0] , \ImageBuffer[3][7] ,
         \ImageBuffer[3][6] , \ImageBuffer[3][5] , \ImageBuffer[3][4] ,
         \ImageBuffer[3][3] , \ImageBuffer[3][2] , \ImageBuffer[3][1] ,
         \ImageBuffer[3][0] , \ImageBuffer[2][7] , \ImageBuffer[2][6] ,
         \ImageBuffer[2][5] , \ImageBuffer[2][4] , \ImageBuffer[2][3] ,
         \ImageBuffer[2][2] , \ImageBuffer[2][1] , \ImageBuffer[2][0] ,
         \ImageBuffer[1][7] , \ImageBuffer[1][6] , \ImageBuffer[1][5] ,
         \ImageBuffer[1][4] , \ImageBuffer[1][3] , \ImageBuffer[1][2] ,
         \ImageBuffer[1][1] , \ImageBuffer[1][0] , \ImageBuffer[0][7] ,
         \ImageBuffer[0][6] , \ImageBuffer[0][5] , \ImageBuffer[0][4] ,
         \ImageBuffer[0][3] , \ImageBuffer[0][2] , \ImageBuffer[0][1] ,
         \ImageBuffer[0][0] , N2673, N2674, N2675, N2695, N2696, N2697, N2701,
         N2702, N2703, N2706, N2707, N2708, N2742, N2743, N2744, N2745, N2746,
         N2747, N2748, N2749, N2750, N2751, N2752, N2753, N2754, N2755, N2756,
         N2757, N2758, N2759, N2760, N2761, N2762, N2763, N2764, N2765, N2766,
         N2767, N2768, N2769, N2770, N2771, N2772, N2773, N2774, N2775, N2776,
         N2777, N2778, N2779, N2780, N2781, N2786, N13064, N13065, N13066,
         N13067, N13068, N13069, N13070, N13071, N13653, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
         n3334, n3335, n3336, n3337, n3338, N2740, N2739, N2738, N2737, N2736,
         N2735, N2734, N2733, N2732, \sub_168_aco/carry[5] ,
         \sub_168_aco/carry[4] , \sub_168_aco/carry[3] ,
         \sub_168_aco/carry[2] , \sub_168_aco/carry[1] , \sub_168_aco/B[0] ,
         \add_162_S2_aco/carry[5] , \add_162_S2_aco/carry[4] ,
         \sub_157_S2_aco/carry[5] , \sub_157_S2_aco/carry[4] ,
         \add_134/carry[5] , \add_134/carry[4] , \add_134/carry[3] ,
         \add_134/carry[2] , \add_122/carry[5] , \add_122/carry[4] ,
         \add_122/carry[3] , \add_122/carry[2] , \add_80/carry[2] ,
         \add_80/carry[3] , \add_80/carry[4] , \add_80/carry[5] ,
         \add_79/carry[5] , \r2549/carry[5] , \r2549/carry[4] ,
         \r2549/carry[3] , \r2549/carry[2] , n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
         n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
         n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n8645, n8646,
         n8647, n8648, n8649, n8650, n8651, n3406, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546,
         n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556,
         n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566,
         n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576,
         n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586,
         n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596,
         n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606,
         n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616,
         n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626,
         n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636,
         n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646,
         n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656,
         n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666,
         n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676,
         n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686,
         n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696,
         n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706,
         n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716,
         n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726,
         n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736,
         n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746,
         n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756,
         n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766,
         n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776,
         n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786,
         n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796,
         n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806,
         n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816,
         n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826,
         n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836,
         n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846,
         n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856,
         n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866,
         n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876,
         n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886,
         n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896,
         n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906,
         n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916,
         n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926,
         n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936,
         n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946,
         n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956,
         n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966,
         n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976,
         n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986,
         n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996,
         n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006,
         n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016,
         n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026,
         n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036,
         n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046,
         n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056,
         n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066,
         n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076,
         n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086,
         n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096,
         n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106,
         n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116,
         n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126,
         n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136,
         n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146,
         n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156,
         n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166,
         n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176,
         n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186,
         n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196,
         n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206,
         n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216,
         n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
         n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236,
         n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246,
         n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
         n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
         n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
         n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
         n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
         n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
         n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
         n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326,
         n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336,
         n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346,
         n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356,
         n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366,
         n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376,
         n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386,
         n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396,
         n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
         n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416,
         n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426,
         n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
         n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
         n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
         n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
         n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
         n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
         n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
         n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
         n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
         n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
         n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
         n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
         n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
         n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
         n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
         n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
         n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
         n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816,
         n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826,
         n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
         n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
         n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
         n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
         n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
         n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
         n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896,
         n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906,
         n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916,
         n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926,
         n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936,
         n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4945, n4946, n4947,
         n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
         n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967,
         n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
         n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
         n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
         n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
         n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
         n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
         n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037,
         n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047,
         n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057,
         n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067,
         n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077,
         n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087,
         n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
         n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107,
         n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117,
         n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127,
         n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137,
         n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147,
         n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157,
         n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167,
         n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
         n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
         n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
         n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207,
         n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217,
         n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227,
         n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237,
         n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247,
         n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257,
         n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267,
         n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277,
         n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287,
         n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297,
         n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307,
         n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317,
         n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327,
         n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337,
         n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347,
         n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357,
         n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367,
         n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377,
         n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387,
         n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397,
         n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407,
         n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417,
         n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427,
         n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437,
         n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447,
         n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457,
         n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467,
         n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477,
         n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487,
         n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497,
         n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507,
         n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517,
         n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527,
         n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537,
         n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547,
         n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557,
         n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567,
         n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577,
         n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587,
         n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597,
         n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607,
         n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617,
         n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627,
         n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637,
         n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647,
         n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657,
         n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667,
         n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677,
         n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687,
         n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697,
         n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707,
         n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717,
         n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727,
         n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737,
         n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747,
         n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757,
         n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767,
         n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777,
         n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787,
         n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797,
         n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807,
         n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817,
         n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827,
         n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837,
         n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847,
         n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857,
         n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867,
         n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877,
         n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887,
         n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897,
         n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907,
         n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917,
         n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927,
         n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937,
         n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947,
         n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957,
         n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967,
         n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977,
         n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987,
         n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997,
         n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007,
         n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017,
         n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027,
         n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037,
         n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047,
         n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057,
         n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067,
         n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077,
         n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087,
         n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097,
         n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107,
         n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117,
         n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127,
         n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137,
         n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147,
         n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157,
         n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167,
         n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177,
         n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187,
         n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197,
         n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207,
         n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217,
         n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227,
         n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237,
         n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247,
         n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257,
         n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267,
         n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277,
         n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287,
         n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297,
         n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307,
         n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317,
         n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327,
         n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337,
         n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347,
         n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357,
         n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367,
         n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377,
         n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387,
         n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397,
         n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407,
         n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417,
         n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427,
         n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437,
         n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447,
         n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457,
         n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467,
         n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477,
         n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487,
         n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497,
         n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507,
         n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517,
         n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527,
         n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537,
         n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547,
         n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557,
         n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
         n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
         n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587,
         n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597,
         n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607,
         n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617,
         n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
         n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
         n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
         n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
         n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
         n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
         n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
         n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
         n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
         n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
         n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
         n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
         n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
         n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
         n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
         n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
         n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
         n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
         n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
         n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
         n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987,
         n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997,
         n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
         n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017,
         n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
         n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037,
         n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047,
         n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
         n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067,
         n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077,
         n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087,
         n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097,
         n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
         n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117,
         n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127,
         n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137,
         n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147,
         n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157,
         n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167,
         n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177,
         n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187,
         n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197,
         n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207,
         n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217,
         n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227,
         n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237,
         n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247,
         n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257,
         n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267,
         n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277,
         n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287,
         n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297,
         n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307,
         n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317,
         n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327,
         n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337,
         n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347,
         n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357,
         n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367,
         n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377,
         n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387,
         n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397,
         n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407,
         n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417,
         n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427,
         n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437,
         n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447,
         n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457,
         n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467,
         n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477,
         n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487,
         n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497,
         n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507,
         n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517,
         n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527,
         n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537,
         n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547,
         n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557,
         n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567,
         n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577,
         n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587,
         n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597,
         n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607,
         n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617,
         n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627,
         n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637,
         n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647,
         n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657,
         n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667,
         n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677,
         n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687,
         n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697,
         n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707,
         n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717,
         n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727,
         n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737,
         n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747,
         n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757,
         n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767,
         n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777,
         n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787,
         n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797,
         n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807,
         n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817,
         n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827,
         n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837,
         n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847,
         n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857,
         n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867,
         n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877,
         n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887,
         n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897,
         n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907,
         n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917,
         n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927,
         n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937,
         n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947,
         n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957,
         n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967,
         n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977,
         n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987,
         n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997,
         n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007,
         n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017,
         n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027,
         n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037,
         n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047,
         n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057,
         n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067,
         n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077,
         n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087,
         n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097,
         n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107,
         n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117,
         n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127,
         n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137,
         n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147,
         n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157,
         n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167,
         n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177,
         n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187,
         n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197,
         n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207,
         n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217,
         n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227,
         n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237,
         n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247,
         n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257,
         n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267,
         n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277,
         n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287,
         n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297,
         n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307,
         n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317,
         n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327,
         n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337,
         n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347,
         n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357,
         n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367,
         n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377,
         n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387,
         n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397,
         n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407,
         n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417,
         n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427,
         n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437,
         n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447,
         n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457,
         n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467,
         n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477,
         n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487,
         n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497,
         n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507,
         n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517,
         n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527,
         n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537,
         n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547,
         n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557,
         n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567,
         n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577,
         n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587,
         n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597,
         n8598, n8599, n8600, n8601, n8602, n8604, n8605, n8606, n8607, n8608,
         n8609, n8610, n8611, n8612, n8613, n8631, n8633, n8635, n8637, n8639,
         n8641, n8643;
  wire   [1:0] state_ns;
  wire   [9:2] sum;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2;
  assign IROM_rd = N2538;

  ADDHX4 \r2549/U1_1_4  ( .A(n5125), .B(\r2549/carry[4] ), .CO(
        \r2549/carry[5] ), .S(N2491) );
  DFFQX1 \counter_reg[1]  ( .D(n3331), .CK(clk), .Q(N2518) );
  DFFQX1 \counter_reg[2]  ( .D(n3330), .CK(clk), .Q(N2519) );
  DFFQX1 \counter_reg[3]  ( .D(n3329), .CK(clk), .Q(N2520) );
  DFFQX1 \counter_reg[0]  ( .D(n3332), .CK(clk), .Q(N2517) );
  DFFQX4 \counter_reg[5]  ( .D(n3327), .CK(clk), .Q(N2522) );
  DFFQX2 \ImageBuffer_reg[61][7]  ( .D(n8092), .CK(clk), .Q(
        \ImageBuffer[61][7] ) );
  DFFQX2 \ImageBuffer_reg[61][6]  ( .D(n8156), .CK(clk), .Q(
        \ImageBuffer[61][6] ) );
  DFFQX2 \ImageBuffer_reg[61][5]  ( .D(n8220), .CK(clk), .Q(
        \ImageBuffer[61][5] ) );
  DFFQX2 \ImageBuffer_reg[61][4]  ( .D(n8284), .CK(clk), .Q(
        \ImageBuffer[61][4] ) );
  DFFQX2 \ImageBuffer_reg[61][3]  ( .D(n8348), .CK(clk), .Q(
        \ImageBuffer[61][3] ) );
  DFFQX2 \ImageBuffer_reg[61][1]  ( .D(n8476), .CK(clk), .Q(
        \ImageBuffer[61][1] ) );
  DFFQX2 \ImageBuffer_reg[57][7]  ( .D(n8096), .CK(clk), .Q(
        \ImageBuffer[57][7] ) );
  DFFQX2 \ImageBuffer_reg[57][6]  ( .D(n8160), .CK(clk), .Q(
        \ImageBuffer[57][6] ) );
  DFFQX2 \ImageBuffer_reg[57][5]  ( .D(n8224), .CK(clk), .Q(
        \ImageBuffer[57][5] ) );
  DFFQX2 \ImageBuffer_reg[57][4]  ( .D(n8288), .CK(clk), .Q(
        \ImageBuffer[57][4] ) );
  DFFQX2 \ImageBuffer_reg[57][3]  ( .D(n8352), .CK(clk), .Q(
        \ImageBuffer[57][3] ) );
  DFFQX2 \ImageBuffer_reg[57][1]  ( .D(n8480), .CK(clk), .Q(
        \ImageBuffer[57][1] ) );
  DFFQX2 \ImageBuffer_reg[53][7]  ( .D(n8100), .CK(clk), .Q(
        \ImageBuffer[53][7] ) );
  DFFQX2 \ImageBuffer_reg[53][6]  ( .D(n8164), .CK(clk), .Q(
        \ImageBuffer[53][6] ) );
  DFFQX2 \ImageBuffer_reg[53][5]  ( .D(n8228), .CK(clk), .Q(
        \ImageBuffer[53][5] ) );
  DFFQX2 \ImageBuffer_reg[53][4]  ( .D(n8292), .CK(clk), .Q(
        \ImageBuffer[53][4] ) );
  DFFQX2 \ImageBuffer_reg[53][3]  ( .D(n8356), .CK(clk), .Q(
        \ImageBuffer[53][3] ) );
  DFFQX2 \ImageBuffer_reg[53][1]  ( .D(n8484), .CK(clk), .Q(
        \ImageBuffer[53][1] ) );
  DFFQX2 \ImageBuffer_reg[49][7]  ( .D(n8104), .CK(clk), .Q(
        \ImageBuffer[49][7] ) );
  DFFQX2 \ImageBuffer_reg[49][6]  ( .D(n8168), .CK(clk), .Q(
        \ImageBuffer[49][6] ) );
  DFFQX2 \ImageBuffer_reg[49][5]  ( .D(n8232), .CK(clk), .Q(
        \ImageBuffer[49][5] ) );
  DFFQX2 \ImageBuffer_reg[49][4]  ( .D(n8296), .CK(clk), .Q(
        \ImageBuffer[49][4] ) );
  DFFQX2 \ImageBuffer_reg[49][3]  ( .D(n8360), .CK(clk), .Q(
        \ImageBuffer[49][3] ) );
  DFFQX2 \ImageBuffer_reg[49][1]  ( .D(n8488), .CK(clk), .Q(
        \ImageBuffer[49][1] ) );
  DFFQX2 \ImageBuffer_reg[45][7]  ( .D(n8108), .CK(clk), .Q(
        \ImageBuffer[45][7] ) );
  DFFQX2 \ImageBuffer_reg[45][6]  ( .D(n8172), .CK(clk), .Q(
        \ImageBuffer[45][6] ) );
  DFFQX2 \ImageBuffer_reg[45][5]  ( .D(n8236), .CK(clk), .Q(
        \ImageBuffer[45][5] ) );
  DFFQX2 \ImageBuffer_reg[45][4]  ( .D(n8300), .CK(clk), .Q(
        \ImageBuffer[45][4] ) );
  DFFQX2 \ImageBuffer_reg[45][3]  ( .D(n8364), .CK(clk), .Q(
        \ImageBuffer[45][3] ) );
  DFFQX2 \ImageBuffer_reg[45][1]  ( .D(n8492), .CK(clk), .Q(
        \ImageBuffer[45][1] ) );
  DFFQX2 \ImageBuffer_reg[41][7]  ( .D(n8112), .CK(clk), .Q(
        \ImageBuffer[41][7] ) );
  DFFQX2 \ImageBuffer_reg[41][6]  ( .D(n8176), .CK(clk), .Q(
        \ImageBuffer[41][6] ) );
  DFFQX2 \ImageBuffer_reg[41][5]  ( .D(n8240), .CK(clk), .Q(
        \ImageBuffer[41][5] ) );
  DFFQX2 \ImageBuffer_reg[41][4]  ( .D(n8304), .CK(clk), .Q(
        \ImageBuffer[41][4] ) );
  DFFQX2 \ImageBuffer_reg[41][3]  ( .D(n8368), .CK(clk), .Q(
        \ImageBuffer[41][3] ) );
  DFFQX2 \ImageBuffer_reg[41][1]  ( .D(n8496), .CK(clk), .Q(
        \ImageBuffer[41][1] ) );
  DFFQX2 \ImageBuffer_reg[37][7]  ( .D(n8116), .CK(clk), .Q(
        \ImageBuffer[37][7] ) );
  DFFQX2 \ImageBuffer_reg[37][6]  ( .D(n8180), .CK(clk), .Q(
        \ImageBuffer[37][6] ) );
  DFFQX2 \ImageBuffer_reg[37][5]  ( .D(n8244), .CK(clk), .Q(
        \ImageBuffer[37][5] ) );
  DFFQX2 \ImageBuffer_reg[37][4]  ( .D(n8308), .CK(clk), .Q(
        \ImageBuffer[37][4] ) );
  DFFQX2 \ImageBuffer_reg[37][3]  ( .D(n8372), .CK(clk), .Q(
        \ImageBuffer[37][3] ) );
  DFFQX2 \ImageBuffer_reg[37][1]  ( .D(n8500), .CK(clk), .Q(
        \ImageBuffer[37][1] ) );
  DFFQX2 \ImageBuffer_reg[33][7]  ( .D(n8120), .CK(clk), .Q(
        \ImageBuffer[33][7] ) );
  DFFQX2 \ImageBuffer_reg[33][6]  ( .D(n8184), .CK(clk), .Q(
        \ImageBuffer[33][6] ) );
  DFFQX2 \ImageBuffer_reg[33][5]  ( .D(n8248), .CK(clk), .Q(
        \ImageBuffer[33][5] ) );
  DFFQX2 \ImageBuffer_reg[33][4]  ( .D(n8312), .CK(clk), .Q(
        \ImageBuffer[33][4] ) );
  DFFQX2 \ImageBuffer_reg[33][3]  ( .D(n8376), .CK(clk), .Q(
        \ImageBuffer[33][3] ) );
  DFFQX2 \ImageBuffer_reg[33][1]  ( .D(n8504), .CK(clk), .Q(
        \ImageBuffer[33][1] ) );
  DFFQX2 \ImageBuffer_reg[29][7]  ( .D(n8124), .CK(clk), .Q(
        \ImageBuffer[29][7] ) );
  DFFQX2 \ImageBuffer_reg[29][6]  ( .D(n8188), .CK(clk), .Q(
        \ImageBuffer[29][6] ) );
  DFFQX2 \ImageBuffer_reg[29][5]  ( .D(n8252), .CK(clk), .Q(
        \ImageBuffer[29][5] ) );
  DFFQX2 \ImageBuffer_reg[29][4]  ( .D(n8316), .CK(clk), .Q(
        \ImageBuffer[29][4] ) );
  DFFQX2 \ImageBuffer_reg[29][3]  ( .D(n8380), .CK(clk), .Q(
        \ImageBuffer[29][3] ) );
  DFFQX2 \ImageBuffer_reg[29][1]  ( .D(n8508), .CK(clk), .Q(
        \ImageBuffer[29][1] ) );
  DFFQX2 \ImageBuffer_reg[25][7]  ( .D(n8128), .CK(clk), .Q(
        \ImageBuffer[25][7] ) );
  DFFQX2 \ImageBuffer_reg[25][6]  ( .D(n8192), .CK(clk), .Q(
        \ImageBuffer[25][6] ) );
  DFFQX2 \ImageBuffer_reg[25][5]  ( .D(n8256), .CK(clk), .Q(
        \ImageBuffer[25][5] ) );
  DFFQX2 \ImageBuffer_reg[25][4]  ( .D(n8320), .CK(clk), .Q(
        \ImageBuffer[25][4] ) );
  DFFQX2 \ImageBuffer_reg[25][3]  ( .D(n8384), .CK(clk), .Q(
        \ImageBuffer[25][3] ) );
  DFFQX2 \ImageBuffer_reg[25][1]  ( .D(n8512), .CK(clk), .Q(
        \ImageBuffer[25][1] ) );
  DFFQX2 \ImageBuffer_reg[21][7]  ( .D(n8132), .CK(clk), .Q(
        \ImageBuffer[21][7] ) );
  DFFQX2 \ImageBuffer_reg[21][6]  ( .D(n8196), .CK(clk), .Q(
        \ImageBuffer[21][6] ) );
  DFFQX2 \ImageBuffer_reg[21][5]  ( .D(n8260), .CK(clk), .Q(
        \ImageBuffer[21][5] ) );
  DFFQX2 \ImageBuffer_reg[21][4]  ( .D(n8324), .CK(clk), .Q(
        \ImageBuffer[21][4] ) );
  DFFQX2 \ImageBuffer_reg[21][3]  ( .D(n8388), .CK(clk), .Q(
        \ImageBuffer[21][3] ) );
  DFFQX2 \ImageBuffer_reg[21][1]  ( .D(n8516), .CK(clk), .Q(
        \ImageBuffer[21][1] ) );
  DFFQX2 \ImageBuffer_reg[17][7]  ( .D(n8136), .CK(clk), .Q(
        \ImageBuffer[17][7] ) );
  DFFQX2 \ImageBuffer_reg[17][6]  ( .D(n8200), .CK(clk), .Q(
        \ImageBuffer[17][6] ) );
  DFFQX2 \ImageBuffer_reg[17][5]  ( .D(n8264), .CK(clk), .Q(
        \ImageBuffer[17][5] ) );
  DFFQX2 \ImageBuffer_reg[17][4]  ( .D(n8328), .CK(clk), .Q(
        \ImageBuffer[17][4] ) );
  DFFQX2 \ImageBuffer_reg[17][3]  ( .D(n8392), .CK(clk), .Q(
        \ImageBuffer[17][3] ) );
  DFFQX2 \ImageBuffer_reg[17][1]  ( .D(n8520), .CK(clk), .Q(
        \ImageBuffer[17][1] ) );
  DFFQX2 \ImageBuffer_reg[13][7]  ( .D(n8140), .CK(clk), .Q(
        \ImageBuffer[13][7] ) );
  DFFQX2 \ImageBuffer_reg[13][6]  ( .D(n8204), .CK(clk), .Q(
        \ImageBuffer[13][6] ) );
  DFFQX2 \ImageBuffer_reg[13][5]  ( .D(n8268), .CK(clk), .Q(
        \ImageBuffer[13][5] ) );
  DFFQX2 \ImageBuffer_reg[13][4]  ( .D(n8332), .CK(clk), .Q(
        \ImageBuffer[13][4] ) );
  DFFQX2 \ImageBuffer_reg[13][3]  ( .D(n8396), .CK(clk), .Q(
        \ImageBuffer[13][3] ) );
  DFFQX2 \ImageBuffer_reg[13][1]  ( .D(n8524), .CK(clk), .Q(
        \ImageBuffer[13][1] ) );
  DFFQX2 \ImageBuffer_reg[9][7]  ( .D(n8144), .CK(clk), .Q(\ImageBuffer[9][7] ) );
  DFFQX2 \ImageBuffer_reg[9][6]  ( .D(n8208), .CK(clk), .Q(\ImageBuffer[9][6] ) );
  DFFQX2 \ImageBuffer_reg[9][5]  ( .D(n8272), .CK(clk), .Q(\ImageBuffer[9][5] ) );
  DFFQX2 \ImageBuffer_reg[9][4]  ( .D(n8336), .CK(clk), .Q(\ImageBuffer[9][4] ) );
  DFFQX2 \ImageBuffer_reg[9][3]  ( .D(n8400), .CK(clk), .Q(\ImageBuffer[9][3] ) );
  DFFQX2 \ImageBuffer_reg[9][1]  ( .D(n8528), .CK(clk), .Q(\ImageBuffer[9][1] ) );
  DFFQX2 \ImageBuffer_reg[5][7]  ( .D(n8148), .CK(clk), .Q(\ImageBuffer[5][7] ) );
  DFFQX2 \ImageBuffer_reg[5][6]  ( .D(n8212), .CK(clk), .Q(\ImageBuffer[5][6] ) );
  DFFQX2 \ImageBuffer_reg[5][5]  ( .D(n8276), .CK(clk), .Q(\ImageBuffer[5][5] ) );
  DFFQX2 \ImageBuffer_reg[5][4]  ( .D(n8340), .CK(clk), .Q(\ImageBuffer[5][4] ) );
  DFFQX2 \ImageBuffer_reg[5][3]  ( .D(n8404), .CK(clk), .Q(\ImageBuffer[5][3] ) );
  DFFQX2 \ImageBuffer_reg[5][1]  ( .D(n8532), .CK(clk), .Q(\ImageBuffer[5][1] ) );
  DFFQX2 \ImageBuffer_reg[1][7]  ( .D(n8152), .CK(clk), .Q(\ImageBuffer[1][7] ) );
  DFFQX2 \ImageBuffer_reg[1][6]  ( .D(n8216), .CK(clk), .Q(\ImageBuffer[1][6] ) );
  DFFQX2 \ImageBuffer_reg[1][5]  ( .D(n8280), .CK(clk), .Q(\ImageBuffer[1][5] ) );
  DFFQX2 \ImageBuffer_reg[1][4]  ( .D(n8344), .CK(clk), .Q(\ImageBuffer[1][4] ) );
  DFFQX2 \ImageBuffer_reg[1][3]  ( .D(n8408), .CK(clk), .Q(\ImageBuffer[1][3] ) );
  DFFQX2 \ImageBuffer_reg[1][1]  ( .D(n8536), .CK(clk), .Q(\ImageBuffer[1][1] ) );
  DFFQX2 \ImageBuffer_reg[63][7]  ( .D(n8090), .CK(clk), .Q(
        \ImageBuffer[63][7] ) );
  DFFQX2 \ImageBuffer_reg[63][6]  ( .D(n8154), .CK(clk), .Q(
        \ImageBuffer[63][6] ) );
  DFFQX2 \ImageBuffer_reg[63][5]  ( .D(n8218), .CK(clk), .Q(
        \ImageBuffer[63][5] ) );
  DFFQX2 \ImageBuffer_reg[63][4]  ( .D(n8282), .CK(clk), .Q(
        \ImageBuffer[63][4] ) );
  DFFQX2 \ImageBuffer_reg[63][3]  ( .D(n8346), .CK(clk), .Q(
        \ImageBuffer[63][3] ) );
  DFFQX2 \ImageBuffer_reg[63][1]  ( .D(n8474), .CK(clk), .Q(
        \ImageBuffer[63][1] ) );
  DFFQX2 \ImageBuffer_reg[59][7]  ( .D(n8094), .CK(clk), .Q(
        \ImageBuffer[59][7] ) );
  DFFQX2 \ImageBuffer_reg[59][6]  ( .D(n8158), .CK(clk), .Q(
        \ImageBuffer[59][6] ) );
  DFFQX2 \ImageBuffer_reg[59][5]  ( .D(n8222), .CK(clk), .Q(
        \ImageBuffer[59][5] ) );
  DFFQX2 \ImageBuffer_reg[59][4]  ( .D(n8286), .CK(clk), .Q(
        \ImageBuffer[59][4] ) );
  DFFQX2 \ImageBuffer_reg[59][3]  ( .D(n8350), .CK(clk), .Q(
        \ImageBuffer[59][3] ) );
  DFFQX2 \ImageBuffer_reg[59][1]  ( .D(n8478), .CK(clk), .Q(
        \ImageBuffer[59][1] ) );
  DFFQX2 \ImageBuffer_reg[55][7]  ( .D(n8098), .CK(clk), .Q(
        \ImageBuffer[55][7] ) );
  DFFQX2 \ImageBuffer_reg[55][6]  ( .D(n8162), .CK(clk), .Q(
        \ImageBuffer[55][6] ) );
  DFFQX2 \ImageBuffer_reg[55][5]  ( .D(n8226), .CK(clk), .Q(
        \ImageBuffer[55][5] ) );
  DFFQX2 \ImageBuffer_reg[55][4]  ( .D(n8290), .CK(clk), .Q(
        \ImageBuffer[55][4] ) );
  DFFQX2 \ImageBuffer_reg[55][3]  ( .D(n8354), .CK(clk), .Q(
        \ImageBuffer[55][3] ) );
  DFFQX2 \ImageBuffer_reg[55][1]  ( .D(n8482), .CK(clk), .Q(
        \ImageBuffer[55][1] ) );
  DFFQX2 \ImageBuffer_reg[51][7]  ( .D(n8102), .CK(clk), .Q(
        \ImageBuffer[51][7] ) );
  DFFQX2 \ImageBuffer_reg[51][6]  ( .D(n8166), .CK(clk), .Q(
        \ImageBuffer[51][6] ) );
  DFFQX2 \ImageBuffer_reg[51][5]  ( .D(n8230), .CK(clk), .Q(
        \ImageBuffer[51][5] ) );
  DFFQX2 \ImageBuffer_reg[51][4]  ( .D(n8294), .CK(clk), .Q(
        \ImageBuffer[51][4] ) );
  DFFQX2 \ImageBuffer_reg[51][3]  ( .D(n8358), .CK(clk), .Q(
        \ImageBuffer[51][3] ) );
  DFFQX2 \ImageBuffer_reg[51][1]  ( .D(n8486), .CK(clk), .Q(
        \ImageBuffer[51][1] ) );
  DFFQX2 \ImageBuffer_reg[47][7]  ( .D(n8106), .CK(clk), .Q(
        \ImageBuffer[47][7] ) );
  DFFQX2 \ImageBuffer_reg[47][6]  ( .D(n8170), .CK(clk), .Q(
        \ImageBuffer[47][6] ) );
  DFFQX2 \ImageBuffer_reg[47][5]  ( .D(n8234), .CK(clk), .Q(
        \ImageBuffer[47][5] ) );
  DFFQX2 \ImageBuffer_reg[47][4]  ( .D(n8298), .CK(clk), .Q(
        \ImageBuffer[47][4] ) );
  DFFQX2 \ImageBuffer_reg[47][3]  ( .D(n8362), .CK(clk), .Q(
        \ImageBuffer[47][3] ) );
  DFFQX2 \ImageBuffer_reg[47][1]  ( .D(n8490), .CK(clk), .Q(
        \ImageBuffer[47][1] ) );
  DFFQX2 \ImageBuffer_reg[43][7]  ( .D(n8110), .CK(clk), .Q(
        \ImageBuffer[43][7] ) );
  DFFQX2 \ImageBuffer_reg[43][6]  ( .D(n8174), .CK(clk), .Q(
        \ImageBuffer[43][6] ) );
  DFFQX2 \ImageBuffer_reg[43][5]  ( .D(n8238), .CK(clk), .Q(
        \ImageBuffer[43][5] ) );
  DFFQX2 \ImageBuffer_reg[43][4]  ( .D(n8302), .CK(clk), .Q(
        \ImageBuffer[43][4] ) );
  DFFQX2 \ImageBuffer_reg[43][3]  ( .D(n8366), .CK(clk), .Q(
        \ImageBuffer[43][3] ) );
  DFFQX2 \ImageBuffer_reg[43][1]  ( .D(n8494), .CK(clk), .Q(
        \ImageBuffer[43][1] ) );
  DFFQX2 \ImageBuffer_reg[39][7]  ( .D(n8114), .CK(clk), .Q(
        \ImageBuffer[39][7] ) );
  DFFQX2 \ImageBuffer_reg[39][6]  ( .D(n8178), .CK(clk), .Q(
        \ImageBuffer[39][6] ) );
  DFFQX2 \ImageBuffer_reg[39][5]  ( .D(n8242), .CK(clk), .Q(
        \ImageBuffer[39][5] ) );
  DFFQX2 \ImageBuffer_reg[39][4]  ( .D(n8306), .CK(clk), .Q(
        \ImageBuffer[39][4] ) );
  DFFQX2 \ImageBuffer_reg[39][3]  ( .D(n8370), .CK(clk), .Q(
        \ImageBuffer[39][3] ) );
  DFFQX2 \ImageBuffer_reg[39][1]  ( .D(n8498), .CK(clk), .Q(
        \ImageBuffer[39][1] ) );
  DFFQX2 \ImageBuffer_reg[35][7]  ( .D(n8118), .CK(clk), .Q(
        \ImageBuffer[35][7] ) );
  DFFQX2 \ImageBuffer_reg[35][6]  ( .D(n8182), .CK(clk), .Q(
        \ImageBuffer[35][6] ) );
  DFFQX2 \ImageBuffer_reg[35][5]  ( .D(n8246), .CK(clk), .Q(
        \ImageBuffer[35][5] ) );
  DFFQX2 \ImageBuffer_reg[35][4]  ( .D(n8310), .CK(clk), .Q(
        \ImageBuffer[35][4] ) );
  DFFQX2 \ImageBuffer_reg[35][3]  ( .D(n8374), .CK(clk), .Q(
        \ImageBuffer[35][3] ) );
  DFFQX2 \ImageBuffer_reg[35][1]  ( .D(n8502), .CK(clk), .Q(
        \ImageBuffer[35][1] ) );
  DFFQX2 \ImageBuffer_reg[31][7]  ( .D(n8122), .CK(clk), .Q(
        \ImageBuffer[31][7] ) );
  DFFQX2 \ImageBuffer_reg[31][6]  ( .D(n8186), .CK(clk), .Q(
        \ImageBuffer[31][6] ) );
  DFFQX2 \ImageBuffer_reg[31][5]  ( .D(n8250), .CK(clk), .Q(
        \ImageBuffer[31][5] ) );
  DFFQX2 \ImageBuffer_reg[31][4]  ( .D(n8314), .CK(clk), .Q(
        \ImageBuffer[31][4] ) );
  DFFQX2 \ImageBuffer_reg[31][3]  ( .D(n8378), .CK(clk), .Q(
        \ImageBuffer[31][3] ) );
  DFFQX2 \ImageBuffer_reg[31][1]  ( .D(n8506), .CK(clk), .Q(
        \ImageBuffer[31][1] ) );
  DFFQX2 \ImageBuffer_reg[27][7]  ( .D(n8126), .CK(clk), .Q(
        \ImageBuffer[27][7] ) );
  DFFQX2 \ImageBuffer_reg[27][6]  ( .D(n8190), .CK(clk), .Q(
        \ImageBuffer[27][6] ) );
  DFFQX2 \ImageBuffer_reg[27][5]  ( .D(n8254), .CK(clk), .Q(
        \ImageBuffer[27][5] ) );
  DFFQX2 \ImageBuffer_reg[27][4]  ( .D(n8318), .CK(clk), .Q(
        \ImageBuffer[27][4] ) );
  DFFQX2 \ImageBuffer_reg[27][3]  ( .D(n8382), .CK(clk), .Q(
        \ImageBuffer[27][3] ) );
  DFFQX2 \ImageBuffer_reg[27][1]  ( .D(n8510), .CK(clk), .Q(
        \ImageBuffer[27][1] ) );
  DFFQX2 \ImageBuffer_reg[23][7]  ( .D(n8130), .CK(clk), .Q(
        \ImageBuffer[23][7] ) );
  DFFQX2 \ImageBuffer_reg[23][6]  ( .D(n8194), .CK(clk), .Q(
        \ImageBuffer[23][6] ) );
  DFFQX2 \ImageBuffer_reg[23][5]  ( .D(n8258), .CK(clk), .Q(
        \ImageBuffer[23][5] ) );
  DFFQX2 \ImageBuffer_reg[23][4]  ( .D(n8322), .CK(clk), .Q(
        \ImageBuffer[23][4] ) );
  DFFQX2 \ImageBuffer_reg[23][3]  ( .D(n8386), .CK(clk), .Q(
        \ImageBuffer[23][3] ) );
  DFFQX2 \ImageBuffer_reg[23][1]  ( .D(n8514), .CK(clk), .Q(
        \ImageBuffer[23][1] ) );
  DFFQX2 \ImageBuffer_reg[19][7]  ( .D(n8134), .CK(clk), .Q(
        \ImageBuffer[19][7] ) );
  DFFQX2 \ImageBuffer_reg[19][6]  ( .D(n8198), .CK(clk), .Q(
        \ImageBuffer[19][6] ) );
  DFFQX2 \ImageBuffer_reg[19][5]  ( .D(n8262), .CK(clk), .Q(
        \ImageBuffer[19][5] ) );
  DFFQX2 \ImageBuffer_reg[19][4]  ( .D(n8326), .CK(clk), .Q(
        \ImageBuffer[19][4] ) );
  DFFQX2 \ImageBuffer_reg[19][3]  ( .D(n8390), .CK(clk), .Q(
        \ImageBuffer[19][3] ) );
  DFFQX2 \ImageBuffer_reg[19][1]  ( .D(n8518), .CK(clk), .Q(
        \ImageBuffer[19][1] ) );
  DFFQX2 \ImageBuffer_reg[15][7]  ( .D(n8138), .CK(clk), .Q(
        \ImageBuffer[15][7] ) );
  DFFQX2 \ImageBuffer_reg[15][6]  ( .D(n8202), .CK(clk), .Q(
        \ImageBuffer[15][6] ) );
  DFFQX2 \ImageBuffer_reg[15][5]  ( .D(n8266), .CK(clk), .Q(
        \ImageBuffer[15][5] ) );
  DFFQX2 \ImageBuffer_reg[15][4]  ( .D(n8330), .CK(clk), .Q(
        \ImageBuffer[15][4] ) );
  DFFQX2 \ImageBuffer_reg[15][3]  ( .D(n8394), .CK(clk), .Q(
        \ImageBuffer[15][3] ) );
  DFFQX2 \ImageBuffer_reg[15][1]  ( .D(n8522), .CK(clk), .Q(
        \ImageBuffer[15][1] ) );
  DFFQX2 \ImageBuffer_reg[11][7]  ( .D(n8142), .CK(clk), .Q(
        \ImageBuffer[11][7] ) );
  DFFQX2 \ImageBuffer_reg[11][6]  ( .D(n8206), .CK(clk), .Q(
        \ImageBuffer[11][6] ) );
  DFFQX2 \ImageBuffer_reg[11][5]  ( .D(n8270), .CK(clk), .Q(
        \ImageBuffer[11][5] ) );
  DFFQX2 \ImageBuffer_reg[11][4]  ( .D(n8334), .CK(clk), .Q(
        \ImageBuffer[11][4] ) );
  DFFQX2 \ImageBuffer_reg[11][3]  ( .D(n8398), .CK(clk), .Q(
        \ImageBuffer[11][3] ) );
  DFFQX2 \ImageBuffer_reg[11][1]  ( .D(n8526), .CK(clk), .Q(
        \ImageBuffer[11][1] ) );
  DFFQX2 \ImageBuffer_reg[7][7]  ( .D(n8146), .CK(clk), .Q(\ImageBuffer[7][7] ) );
  DFFQX2 \ImageBuffer_reg[7][6]  ( .D(n8210), .CK(clk), .Q(\ImageBuffer[7][6] ) );
  DFFQX2 \ImageBuffer_reg[7][5]  ( .D(n8274), .CK(clk), .Q(\ImageBuffer[7][5] ) );
  DFFQX2 \ImageBuffer_reg[7][4]  ( .D(n8338), .CK(clk), .Q(\ImageBuffer[7][4] ) );
  DFFQX2 \ImageBuffer_reg[7][3]  ( .D(n8402), .CK(clk), .Q(\ImageBuffer[7][3] ) );
  DFFQX2 \ImageBuffer_reg[7][1]  ( .D(n8530), .CK(clk), .Q(\ImageBuffer[7][1] ) );
  DFFQX2 \ImageBuffer_reg[3][7]  ( .D(n8150), .CK(clk), .Q(\ImageBuffer[3][7] ) );
  DFFQX2 \ImageBuffer_reg[3][6]  ( .D(n8214), .CK(clk), .Q(\ImageBuffer[3][6] ) );
  DFFQX2 \ImageBuffer_reg[3][5]  ( .D(n8278), .CK(clk), .Q(\ImageBuffer[3][5] ) );
  DFFQX2 \ImageBuffer_reg[3][4]  ( .D(n8342), .CK(clk), .Q(\ImageBuffer[3][4] ) );
  DFFQX2 \ImageBuffer_reg[3][3]  ( .D(n8406), .CK(clk), .Q(\ImageBuffer[3][3] ) );
  DFFQX2 \ImageBuffer_reg[3][1]  ( .D(n8534), .CK(clk), .Q(\ImageBuffer[3][1] ) );
  DFFQX2 \ImageBuffer_reg[60][7]  ( .D(n8093), .CK(clk), .Q(
        \ImageBuffer[60][7] ) );
  DFFQX2 \ImageBuffer_reg[60][6]  ( .D(n8157), .CK(clk), .Q(
        \ImageBuffer[60][6] ) );
  DFFQX2 \ImageBuffer_reg[60][5]  ( .D(n8221), .CK(clk), .Q(
        \ImageBuffer[60][5] ) );
  DFFQX2 \ImageBuffer_reg[60][4]  ( .D(n8285), .CK(clk), .Q(
        \ImageBuffer[60][4] ) );
  DFFQX2 \ImageBuffer_reg[60][3]  ( .D(n8349), .CK(clk), .Q(
        \ImageBuffer[60][3] ) );
  DFFQX2 \ImageBuffer_reg[60][1]  ( .D(n8477), .CK(clk), .Q(
        \ImageBuffer[60][1] ) );
  DFFQX2 \ImageBuffer_reg[56][7]  ( .D(n8097), .CK(clk), .Q(
        \ImageBuffer[56][7] ) );
  DFFQX2 \ImageBuffer_reg[56][6]  ( .D(n8161), .CK(clk), .Q(
        \ImageBuffer[56][6] ) );
  DFFQX2 \ImageBuffer_reg[56][5]  ( .D(n8225), .CK(clk), .Q(
        \ImageBuffer[56][5] ) );
  DFFQX2 \ImageBuffer_reg[56][4]  ( .D(n8289), .CK(clk), .Q(
        \ImageBuffer[56][4] ) );
  DFFQX2 \ImageBuffer_reg[56][3]  ( .D(n8353), .CK(clk), .Q(
        \ImageBuffer[56][3] ) );
  DFFQX2 \ImageBuffer_reg[56][1]  ( .D(n8481), .CK(clk), .Q(
        \ImageBuffer[56][1] ) );
  DFFQX2 \ImageBuffer_reg[52][7]  ( .D(n8101), .CK(clk), .Q(
        \ImageBuffer[52][7] ) );
  DFFQX2 \ImageBuffer_reg[52][6]  ( .D(n8165), .CK(clk), .Q(
        \ImageBuffer[52][6] ) );
  DFFQX2 \ImageBuffer_reg[52][5]  ( .D(n8229), .CK(clk), .Q(
        \ImageBuffer[52][5] ) );
  DFFQX2 \ImageBuffer_reg[52][4]  ( .D(n8293), .CK(clk), .Q(
        \ImageBuffer[52][4] ) );
  DFFQX2 \ImageBuffer_reg[52][3]  ( .D(n8357), .CK(clk), .Q(
        \ImageBuffer[52][3] ) );
  DFFQX2 \ImageBuffer_reg[52][1]  ( .D(n8485), .CK(clk), .Q(
        \ImageBuffer[52][1] ) );
  DFFQX2 \ImageBuffer_reg[48][7]  ( .D(n8105), .CK(clk), .Q(
        \ImageBuffer[48][7] ) );
  DFFQX2 \ImageBuffer_reg[48][6]  ( .D(n8169), .CK(clk), .Q(
        \ImageBuffer[48][6] ) );
  DFFQX2 \ImageBuffer_reg[48][5]  ( .D(n8233), .CK(clk), .Q(
        \ImageBuffer[48][5] ) );
  DFFQX2 \ImageBuffer_reg[48][4]  ( .D(n8297), .CK(clk), .Q(
        \ImageBuffer[48][4] ) );
  DFFQX2 \ImageBuffer_reg[48][3]  ( .D(n8361), .CK(clk), .Q(
        \ImageBuffer[48][3] ) );
  DFFQX2 \ImageBuffer_reg[48][1]  ( .D(n8489), .CK(clk), .Q(
        \ImageBuffer[48][1] ) );
  DFFQX2 \ImageBuffer_reg[44][7]  ( .D(n8109), .CK(clk), .Q(
        \ImageBuffer[44][7] ) );
  DFFQX2 \ImageBuffer_reg[44][6]  ( .D(n8173), .CK(clk), .Q(
        \ImageBuffer[44][6] ) );
  DFFQX2 \ImageBuffer_reg[44][5]  ( .D(n8237), .CK(clk), .Q(
        \ImageBuffer[44][5] ) );
  DFFQX2 \ImageBuffer_reg[44][4]  ( .D(n8301), .CK(clk), .Q(
        \ImageBuffer[44][4] ) );
  DFFQX2 \ImageBuffer_reg[44][3]  ( .D(n8365), .CK(clk), .Q(
        \ImageBuffer[44][3] ) );
  DFFQX2 \ImageBuffer_reg[44][1]  ( .D(n8493), .CK(clk), .Q(
        \ImageBuffer[44][1] ) );
  DFFQX2 \ImageBuffer_reg[40][7]  ( .D(n8113), .CK(clk), .Q(
        \ImageBuffer[40][7] ) );
  DFFQX2 \ImageBuffer_reg[40][6]  ( .D(n8177), .CK(clk), .Q(
        \ImageBuffer[40][6] ) );
  DFFQX2 \ImageBuffer_reg[40][5]  ( .D(n8241), .CK(clk), .Q(
        \ImageBuffer[40][5] ) );
  DFFQX2 \ImageBuffer_reg[40][4]  ( .D(n8305), .CK(clk), .Q(
        \ImageBuffer[40][4] ) );
  DFFQX2 \ImageBuffer_reg[40][3]  ( .D(n8369), .CK(clk), .Q(
        \ImageBuffer[40][3] ) );
  DFFQX2 \ImageBuffer_reg[40][1]  ( .D(n8497), .CK(clk), .Q(
        \ImageBuffer[40][1] ) );
  DFFQX2 \ImageBuffer_reg[36][7]  ( .D(n8117), .CK(clk), .Q(
        \ImageBuffer[36][7] ) );
  DFFQX2 \ImageBuffer_reg[36][6]  ( .D(n8181), .CK(clk), .Q(
        \ImageBuffer[36][6] ) );
  DFFQX2 \ImageBuffer_reg[36][5]  ( .D(n8245), .CK(clk), .Q(
        \ImageBuffer[36][5] ) );
  DFFQX2 \ImageBuffer_reg[36][4]  ( .D(n8309), .CK(clk), .Q(
        \ImageBuffer[36][4] ) );
  DFFQX2 \ImageBuffer_reg[36][3]  ( .D(n8373), .CK(clk), .Q(
        \ImageBuffer[36][3] ) );
  DFFQX2 \ImageBuffer_reg[36][1]  ( .D(n8501), .CK(clk), .Q(
        \ImageBuffer[36][1] ) );
  DFFQX2 \ImageBuffer_reg[32][7]  ( .D(n8121), .CK(clk), .Q(
        \ImageBuffer[32][7] ) );
  DFFQX2 \ImageBuffer_reg[32][6]  ( .D(n8185), .CK(clk), .Q(
        \ImageBuffer[32][6] ) );
  DFFQX2 \ImageBuffer_reg[32][5]  ( .D(n8249), .CK(clk), .Q(
        \ImageBuffer[32][5] ) );
  DFFQX2 \ImageBuffer_reg[32][4]  ( .D(n8313), .CK(clk), .Q(
        \ImageBuffer[32][4] ) );
  DFFQX2 \ImageBuffer_reg[32][3]  ( .D(n8377), .CK(clk), .Q(
        \ImageBuffer[32][3] ) );
  DFFQX2 \ImageBuffer_reg[32][1]  ( .D(n8505), .CK(clk), .Q(
        \ImageBuffer[32][1] ) );
  DFFQX2 \ImageBuffer_reg[28][7]  ( .D(n8125), .CK(clk), .Q(
        \ImageBuffer[28][7] ) );
  DFFQX2 \ImageBuffer_reg[28][6]  ( .D(n8189), .CK(clk), .Q(
        \ImageBuffer[28][6] ) );
  DFFQX2 \ImageBuffer_reg[28][5]  ( .D(n8253), .CK(clk), .Q(
        \ImageBuffer[28][5] ) );
  DFFQX2 \ImageBuffer_reg[28][4]  ( .D(n8317), .CK(clk), .Q(
        \ImageBuffer[28][4] ) );
  DFFQX2 \ImageBuffer_reg[28][3]  ( .D(n8381), .CK(clk), .Q(
        \ImageBuffer[28][3] ) );
  DFFQX2 \ImageBuffer_reg[28][1]  ( .D(n8509), .CK(clk), .Q(
        \ImageBuffer[28][1] ) );
  DFFQX2 \ImageBuffer_reg[24][7]  ( .D(n8129), .CK(clk), .Q(
        \ImageBuffer[24][7] ) );
  DFFQX2 \ImageBuffer_reg[24][6]  ( .D(n8193), .CK(clk), .Q(
        \ImageBuffer[24][6] ) );
  DFFQX2 \ImageBuffer_reg[24][5]  ( .D(n8257), .CK(clk), .Q(
        \ImageBuffer[24][5] ) );
  DFFQX2 \ImageBuffer_reg[24][4]  ( .D(n8321), .CK(clk), .Q(
        \ImageBuffer[24][4] ) );
  DFFQX2 \ImageBuffer_reg[24][3]  ( .D(n8385), .CK(clk), .Q(
        \ImageBuffer[24][3] ) );
  DFFQX2 \ImageBuffer_reg[24][1]  ( .D(n8513), .CK(clk), .Q(
        \ImageBuffer[24][1] ) );
  DFFQX2 \ImageBuffer_reg[20][7]  ( .D(n8133), .CK(clk), .Q(
        \ImageBuffer[20][7] ) );
  DFFQX2 \ImageBuffer_reg[20][6]  ( .D(n8197), .CK(clk), .Q(
        \ImageBuffer[20][6] ) );
  DFFQX2 \ImageBuffer_reg[20][5]  ( .D(n8261), .CK(clk), .Q(
        \ImageBuffer[20][5] ) );
  DFFQX2 \ImageBuffer_reg[20][4]  ( .D(n8325), .CK(clk), .Q(
        \ImageBuffer[20][4] ) );
  DFFQX2 \ImageBuffer_reg[20][3]  ( .D(n8389), .CK(clk), .Q(
        \ImageBuffer[20][3] ) );
  DFFQX2 \ImageBuffer_reg[20][1]  ( .D(n8517), .CK(clk), .Q(
        \ImageBuffer[20][1] ) );
  DFFQX2 \ImageBuffer_reg[16][7]  ( .D(n8137), .CK(clk), .Q(
        \ImageBuffer[16][7] ) );
  DFFQX2 \ImageBuffer_reg[16][6]  ( .D(n8201), .CK(clk), .Q(
        \ImageBuffer[16][6] ) );
  DFFQX2 \ImageBuffer_reg[16][5]  ( .D(n8265), .CK(clk), .Q(
        \ImageBuffer[16][5] ) );
  DFFQX2 \ImageBuffer_reg[16][4]  ( .D(n8329), .CK(clk), .Q(
        \ImageBuffer[16][4] ) );
  DFFQX2 \ImageBuffer_reg[16][3]  ( .D(n8393), .CK(clk), .Q(
        \ImageBuffer[16][3] ) );
  DFFQX2 \ImageBuffer_reg[16][1]  ( .D(n8521), .CK(clk), .Q(
        \ImageBuffer[16][1] ) );
  DFFQX2 \ImageBuffer_reg[12][7]  ( .D(n8141), .CK(clk), .Q(
        \ImageBuffer[12][7] ) );
  DFFQX2 \ImageBuffer_reg[12][6]  ( .D(n8205), .CK(clk), .Q(
        \ImageBuffer[12][6] ) );
  DFFQX2 \ImageBuffer_reg[12][5]  ( .D(n8269), .CK(clk), .Q(
        \ImageBuffer[12][5] ) );
  DFFQX2 \ImageBuffer_reg[12][4]  ( .D(n8333), .CK(clk), .Q(
        \ImageBuffer[12][4] ) );
  DFFQX2 \ImageBuffer_reg[12][3]  ( .D(n8397), .CK(clk), .Q(
        \ImageBuffer[12][3] ) );
  DFFQX2 \ImageBuffer_reg[12][1]  ( .D(n8525), .CK(clk), .Q(
        \ImageBuffer[12][1] ) );
  DFFQX2 \ImageBuffer_reg[8][7]  ( .D(n8145), .CK(clk), .Q(\ImageBuffer[8][7] ) );
  DFFQX2 \ImageBuffer_reg[8][6]  ( .D(n8209), .CK(clk), .Q(\ImageBuffer[8][6] ) );
  DFFQX2 \ImageBuffer_reg[8][5]  ( .D(n8273), .CK(clk), .Q(\ImageBuffer[8][5] ) );
  DFFQX2 \ImageBuffer_reg[8][4]  ( .D(n8337), .CK(clk), .Q(\ImageBuffer[8][4] ) );
  DFFQX2 \ImageBuffer_reg[8][3]  ( .D(n8401), .CK(clk), .Q(\ImageBuffer[8][3] ) );
  DFFQX2 \ImageBuffer_reg[8][1]  ( .D(n8529), .CK(clk), .Q(\ImageBuffer[8][1] ) );
  DFFQX2 \ImageBuffer_reg[4][7]  ( .D(n8149), .CK(clk), .Q(\ImageBuffer[4][7] ) );
  DFFQX2 \ImageBuffer_reg[4][6]  ( .D(n8213), .CK(clk), .Q(\ImageBuffer[4][6] ) );
  DFFQX2 \ImageBuffer_reg[4][5]  ( .D(n8277), .CK(clk), .Q(\ImageBuffer[4][5] ) );
  DFFQX2 \ImageBuffer_reg[4][4]  ( .D(n8341), .CK(clk), .Q(\ImageBuffer[4][4] ) );
  DFFQX2 \ImageBuffer_reg[4][3]  ( .D(n8405), .CK(clk), .Q(\ImageBuffer[4][3] ) );
  DFFQX2 \ImageBuffer_reg[4][1]  ( .D(n8533), .CK(clk), .Q(\ImageBuffer[4][1] ) );
  DFFQX2 \ImageBuffer_reg[0][7]  ( .D(n8153), .CK(clk), .Q(\ImageBuffer[0][7] ) );
  DFFQX2 \ImageBuffer_reg[0][6]  ( .D(n8217), .CK(clk), .Q(\ImageBuffer[0][6] ) );
  DFFQX2 \ImageBuffer_reg[0][5]  ( .D(n8281), .CK(clk), .Q(\ImageBuffer[0][5] ) );
  DFFQX2 \ImageBuffer_reg[0][4]  ( .D(n8345), .CK(clk), .Q(\ImageBuffer[0][4] ) );
  DFFQX2 \ImageBuffer_reg[0][3]  ( .D(n8409), .CK(clk), .Q(\ImageBuffer[0][3] ) );
  DFFQX2 \ImageBuffer_reg[0][1]  ( .D(n8537), .CK(clk), .Q(\ImageBuffer[0][1] ) );
  DFFQX2 \ImageBuffer_reg[62][7]  ( .D(n8091), .CK(clk), .Q(
        \ImageBuffer[62][7] ) );
  DFFQX2 \ImageBuffer_reg[62][6]  ( .D(n8155), .CK(clk), .Q(
        \ImageBuffer[62][6] ) );
  DFFQX2 \ImageBuffer_reg[62][5]  ( .D(n8219), .CK(clk), .Q(
        \ImageBuffer[62][5] ) );
  DFFQX2 \ImageBuffer_reg[62][4]  ( .D(n8283), .CK(clk), .Q(
        \ImageBuffer[62][4] ) );
  DFFQX2 \ImageBuffer_reg[62][3]  ( .D(n8347), .CK(clk), .Q(
        \ImageBuffer[62][3] ) );
  DFFQX2 \ImageBuffer_reg[62][1]  ( .D(n8475), .CK(clk), .Q(
        \ImageBuffer[62][1] ) );
  DFFQX2 \ImageBuffer_reg[58][7]  ( .D(n8095), .CK(clk), .Q(
        \ImageBuffer[58][7] ) );
  DFFQX2 \ImageBuffer_reg[58][6]  ( .D(n8159), .CK(clk), .Q(
        \ImageBuffer[58][6] ) );
  DFFQX2 \ImageBuffer_reg[58][5]  ( .D(n8223), .CK(clk), .Q(
        \ImageBuffer[58][5] ) );
  DFFQX2 \ImageBuffer_reg[58][4]  ( .D(n8287), .CK(clk), .Q(
        \ImageBuffer[58][4] ) );
  DFFQX2 \ImageBuffer_reg[58][3]  ( .D(n8351), .CK(clk), .Q(
        \ImageBuffer[58][3] ) );
  DFFQX2 \ImageBuffer_reg[58][1]  ( .D(n8479), .CK(clk), .Q(
        \ImageBuffer[58][1] ) );
  DFFQX2 \ImageBuffer_reg[54][7]  ( .D(n8099), .CK(clk), .Q(
        \ImageBuffer[54][7] ) );
  DFFQX2 \ImageBuffer_reg[54][6]  ( .D(n8163), .CK(clk), .Q(
        \ImageBuffer[54][6] ) );
  DFFQX2 \ImageBuffer_reg[54][5]  ( .D(n8227), .CK(clk), .Q(
        \ImageBuffer[54][5] ) );
  DFFQX2 \ImageBuffer_reg[54][4]  ( .D(n8291), .CK(clk), .Q(
        \ImageBuffer[54][4] ) );
  DFFQX2 \ImageBuffer_reg[54][3]  ( .D(n8355), .CK(clk), .Q(
        \ImageBuffer[54][3] ) );
  DFFQX2 \ImageBuffer_reg[54][1]  ( .D(n8483), .CK(clk), .Q(
        \ImageBuffer[54][1] ) );
  DFFQX2 \ImageBuffer_reg[50][7]  ( .D(n8103), .CK(clk), .Q(
        \ImageBuffer[50][7] ) );
  DFFQX2 \ImageBuffer_reg[50][6]  ( .D(n8167), .CK(clk), .Q(
        \ImageBuffer[50][6] ) );
  DFFQX2 \ImageBuffer_reg[50][5]  ( .D(n8231), .CK(clk), .Q(
        \ImageBuffer[50][5] ) );
  DFFQX2 \ImageBuffer_reg[50][4]  ( .D(n8295), .CK(clk), .Q(
        \ImageBuffer[50][4] ) );
  DFFQX2 \ImageBuffer_reg[50][3]  ( .D(n8359), .CK(clk), .Q(
        \ImageBuffer[50][3] ) );
  DFFQX2 \ImageBuffer_reg[50][1]  ( .D(n8487), .CK(clk), .Q(
        \ImageBuffer[50][1] ) );
  DFFQX2 \ImageBuffer_reg[46][7]  ( .D(n8107), .CK(clk), .Q(
        \ImageBuffer[46][7] ) );
  DFFQX2 \ImageBuffer_reg[46][6]  ( .D(n8171), .CK(clk), .Q(
        \ImageBuffer[46][6] ) );
  DFFQX2 \ImageBuffer_reg[46][5]  ( .D(n8235), .CK(clk), .Q(
        \ImageBuffer[46][5] ) );
  DFFQX2 \ImageBuffer_reg[46][4]  ( .D(n8299), .CK(clk), .Q(
        \ImageBuffer[46][4] ) );
  DFFQX2 \ImageBuffer_reg[46][3]  ( .D(n8363), .CK(clk), .Q(
        \ImageBuffer[46][3] ) );
  DFFQX2 \ImageBuffer_reg[46][1]  ( .D(n8491), .CK(clk), .Q(
        \ImageBuffer[46][1] ) );
  DFFQX2 \ImageBuffer_reg[42][7]  ( .D(n8111), .CK(clk), .Q(
        \ImageBuffer[42][7] ) );
  DFFQX2 \ImageBuffer_reg[42][6]  ( .D(n8175), .CK(clk), .Q(
        \ImageBuffer[42][6] ) );
  DFFQX2 \ImageBuffer_reg[42][5]  ( .D(n8239), .CK(clk), .Q(
        \ImageBuffer[42][5] ) );
  DFFQX2 \ImageBuffer_reg[42][4]  ( .D(n8303), .CK(clk), .Q(
        \ImageBuffer[42][4] ) );
  DFFQX2 \ImageBuffer_reg[42][3]  ( .D(n8367), .CK(clk), .Q(
        \ImageBuffer[42][3] ) );
  DFFQX2 \ImageBuffer_reg[42][1]  ( .D(n8495), .CK(clk), .Q(
        \ImageBuffer[42][1] ) );
  DFFQX2 \ImageBuffer_reg[38][6]  ( .D(n8179), .CK(clk), .Q(
        \ImageBuffer[38][6] ) );
  DFFQX2 \ImageBuffer_reg[38][5]  ( .D(n8243), .CK(clk), .Q(
        \ImageBuffer[38][5] ) );
  DFFQX2 \ImageBuffer_reg[38][4]  ( .D(n8307), .CK(clk), .Q(
        \ImageBuffer[38][4] ) );
  DFFQX2 \ImageBuffer_reg[38][3]  ( .D(n8371), .CK(clk), .Q(
        \ImageBuffer[38][3] ) );
  DFFQX2 \ImageBuffer_reg[38][1]  ( .D(n8499), .CK(clk), .Q(
        \ImageBuffer[38][1] ) );
  DFFQX2 \ImageBuffer_reg[34][7]  ( .D(n8119), .CK(clk), .Q(
        \ImageBuffer[34][7] ) );
  DFFQX2 \ImageBuffer_reg[34][6]  ( .D(n8183), .CK(clk), .Q(
        \ImageBuffer[34][6] ) );
  DFFQX2 \ImageBuffer_reg[34][5]  ( .D(n8247), .CK(clk), .Q(
        \ImageBuffer[34][5] ) );
  DFFQX2 \ImageBuffer_reg[34][4]  ( .D(n8311), .CK(clk), .Q(
        \ImageBuffer[34][4] ) );
  DFFQX2 \ImageBuffer_reg[34][3]  ( .D(n8375), .CK(clk), .Q(
        \ImageBuffer[34][3] ) );
  DFFQX2 \ImageBuffer_reg[34][1]  ( .D(n8503), .CK(clk), .Q(
        \ImageBuffer[34][1] ) );
  DFFQX2 \ImageBuffer_reg[30][7]  ( .D(n8123), .CK(clk), .Q(
        \ImageBuffer[30][7] ) );
  DFFQX2 \ImageBuffer_reg[30][6]  ( .D(n8187), .CK(clk), .Q(
        \ImageBuffer[30][6] ) );
  DFFQX2 \ImageBuffer_reg[30][5]  ( .D(n8251), .CK(clk), .Q(
        \ImageBuffer[30][5] ) );
  DFFQX2 \ImageBuffer_reg[30][4]  ( .D(n8315), .CK(clk), .Q(
        \ImageBuffer[30][4] ) );
  DFFQX2 \ImageBuffer_reg[30][3]  ( .D(n8379), .CK(clk), .Q(
        \ImageBuffer[30][3] ) );
  DFFQX2 \ImageBuffer_reg[30][1]  ( .D(n8507), .CK(clk), .Q(
        \ImageBuffer[30][1] ) );
  DFFQX2 \ImageBuffer_reg[26][7]  ( .D(n8127), .CK(clk), .Q(
        \ImageBuffer[26][7] ) );
  DFFQX2 \ImageBuffer_reg[26][6]  ( .D(n8191), .CK(clk), .Q(
        \ImageBuffer[26][6] ) );
  DFFQX2 \ImageBuffer_reg[26][5]  ( .D(n8255), .CK(clk), .Q(
        \ImageBuffer[26][5] ) );
  DFFQX2 \ImageBuffer_reg[26][4]  ( .D(n8319), .CK(clk), .Q(
        \ImageBuffer[26][4] ) );
  DFFQX2 \ImageBuffer_reg[26][3]  ( .D(n8383), .CK(clk), .Q(
        \ImageBuffer[26][3] ) );
  DFFQX2 \ImageBuffer_reg[26][1]  ( .D(n8511), .CK(clk), .Q(
        \ImageBuffer[26][1] ) );
  DFFQX2 \ImageBuffer_reg[22][7]  ( .D(n8131), .CK(clk), .Q(
        \ImageBuffer[22][7] ) );
  DFFQX2 \ImageBuffer_reg[22][6]  ( .D(n8195), .CK(clk), .Q(
        \ImageBuffer[22][6] ) );
  DFFQX2 \ImageBuffer_reg[22][5]  ( .D(n8259), .CK(clk), .Q(
        \ImageBuffer[22][5] ) );
  DFFQX2 \ImageBuffer_reg[22][4]  ( .D(n8323), .CK(clk), .Q(
        \ImageBuffer[22][4] ) );
  DFFQX2 \ImageBuffer_reg[22][3]  ( .D(n8387), .CK(clk), .Q(
        \ImageBuffer[22][3] ) );
  DFFQX2 \ImageBuffer_reg[22][1]  ( .D(n8515), .CK(clk), .Q(
        \ImageBuffer[22][1] ) );
  DFFQX2 \ImageBuffer_reg[18][7]  ( .D(n8135), .CK(clk), .Q(
        \ImageBuffer[18][7] ) );
  DFFQX2 \ImageBuffer_reg[18][6]  ( .D(n8199), .CK(clk), .Q(
        \ImageBuffer[18][6] ) );
  DFFQX2 \ImageBuffer_reg[18][5]  ( .D(n8263), .CK(clk), .Q(
        \ImageBuffer[18][5] ) );
  DFFQX2 \ImageBuffer_reg[18][4]  ( .D(n8327), .CK(clk), .Q(
        \ImageBuffer[18][4] ) );
  DFFQX2 \ImageBuffer_reg[18][3]  ( .D(n8391), .CK(clk), .Q(
        \ImageBuffer[18][3] ) );
  DFFQX2 \ImageBuffer_reg[18][1]  ( .D(n8519), .CK(clk), .Q(
        \ImageBuffer[18][1] ) );
  DFFQX2 \ImageBuffer_reg[14][7]  ( .D(n8139), .CK(clk), .Q(
        \ImageBuffer[14][7] ) );
  DFFQX2 \ImageBuffer_reg[14][6]  ( .D(n8203), .CK(clk), .Q(
        \ImageBuffer[14][6] ) );
  DFFQX2 \ImageBuffer_reg[14][5]  ( .D(n8267), .CK(clk), .Q(
        \ImageBuffer[14][5] ) );
  DFFQX2 \ImageBuffer_reg[14][4]  ( .D(n8331), .CK(clk), .Q(
        \ImageBuffer[14][4] ) );
  DFFQX2 \ImageBuffer_reg[14][3]  ( .D(n8395), .CK(clk), .Q(
        \ImageBuffer[14][3] ) );
  DFFQX2 \ImageBuffer_reg[14][1]  ( .D(n8523), .CK(clk), .Q(
        \ImageBuffer[14][1] ) );
  DFFQX2 \ImageBuffer_reg[10][7]  ( .D(n8143), .CK(clk), .Q(
        \ImageBuffer[10][7] ) );
  DFFQX2 \ImageBuffer_reg[10][6]  ( .D(n8207), .CK(clk), .Q(
        \ImageBuffer[10][6] ) );
  DFFQX2 \ImageBuffer_reg[10][5]  ( .D(n8271), .CK(clk), .Q(
        \ImageBuffer[10][5] ) );
  DFFQX2 \ImageBuffer_reg[10][4]  ( .D(n8335), .CK(clk), .Q(
        \ImageBuffer[10][4] ) );
  DFFQX2 \ImageBuffer_reg[10][3]  ( .D(n8399), .CK(clk), .Q(
        \ImageBuffer[10][3] ) );
  DFFQX2 \ImageBuffer_reg[10][1]  ( .D(n8527), .CK(clk), .Q(
        \ImageBuffer[10][1] ) );
  DFFQX2 \ImageBuffer_reg[6][7]  ( .D(n8147), .CK(clk), .Q(\ImageBuffer[6][7] ) );
  DFFQX2 \ImageBuffer_reg[6][6]  ( .D(n8211), .CK(clk), .Q(\ImageBuffer[6][6] ) );
  DFFQX2 \ImageBuffer_reg[6][5]  ( .D(n8275), .CK(clk), .Q(\ImageBuffer[6][5] ) );
  DFFQX2 \ImageBuffer_reg[6][4]  ( .D(n8339), .CK(clk), .Q(\ImageBuffer[6][4] ) );
  DFFQX2 \ImageBuffer_reg[6][3]  ( .D(n8403), .CK(clk), .Q(\ImageBuffer[6][3] ) );
  DFFQX2 \ImageBuffer_reg[6][1]  ( .D(n8531), .CK(clk), .Q(\ImageBuffer[6][1] ) );
  DFFQX2 \ImageBuffer_reg[2][7]  ( .D(n8151), .CK(clk), .Q(\ImageBuffer[2][7] ) );
  DFFQX2 \ImageBuffer_reg[2][6]  ( .D(n8215), .CK(clk), .Q(\ImageBuffer[2][6] ) );
  DFFQX2 \ImageBuffer_reg[2][5]  ( .D(n8279), .CK(clk), .Q(\ImageBuffer[2][5] ) );
  DFFQX2 \ImageBuffer_reg[2][4]  ( .D(n8343), .CK(clk), .Q(\ImageBuffer[2][4] ) );
  DFFQX2 \ImageBuffer_reg[2][3]  ( .D(n8407), .CK(clk), .Q(\ImageBuffer[2][3] ) );
  DFFQX2 \ImageBuffer_reg[2][1]  ( .D(n8535), .CK(clk), .Q(\ImageBuffer[2][1] ) );
  DFFQX2 \ImageBuffer_reg[61][2]  ( .D(n8412), .CK(clk), .Q(
        \ImageBuffer[61][2] ) );
  DFFQX2 \ImageBuffer_reg[57][2]  ( .D(n8416), .CK(clk), .Q(
        \ImageBuffer[57][2] ) );
  DFFQX2 \ImageBuffer_reg[57][0]  ( .D(n8544), .CK(clk), .Q(
        \ImageBuffer[57][0] ) );
  DFFQX2 \ImageBuffer_reg[53][0]  ( .D(n8548), .CK(clk), .Q(
        \ImageBuffer[53][0] ) );
  DFFQX2 \ImageBuffer_reg[49][2]  ( .D(n8424), .CK(clk), .Q(
        \ImageBuffer[49][2] ) );
  DFFQX2 \ImageBuffer_reg[49][0]  ( .D(n8552), .CK(clk), .Q(
        \ImageBuffer[49][0] ) );
  DFFQX2 \ImageBuffer_reg[45][0]  ( .D(n8556), .CK(clk), .Q(
        \ImageBuffer[45][0] ) );
  DFFQX2 \ImageBuffer_reg[41][0]  ( .D(n8560), .CK(clk), .Q(
        \ImageBuffer[41][0] ) );
  DFFQX2 \ImageBuffer_reg[37][2]  ( .D(n8436), .CK(clk), .Q(
        \ImageBuffer[37][2] ) );
  DFFQX2 \ImageBuffer_reg[37][0]  ( .D(n8564), .CK(clk), .Q(
        \ImageBuffer[37][0] ) );
  DFFQX2 \ImageBuffer_reg[33][0]  ( .D(n8568), .CK(clk), .Q(
        \ImageBuffer[33][0] ) );
  DFFQX2 \ImageBuffer_reg[29][0]  ( .D(n8572), .CK(clk), .Q(
        \ImageBuffer[29][0] ) );
  DFFQX2 \ImageBuffer_reg[25][2]  ( .D(n8448), .CK(clk), .Q(
        \ImageBuffer[25][2] ) );
  DFFQX2 \ImageBuffer_reg[25][0]  ( .D(n8576), .CK(clk), .Q(
        \ImageBuffer[25][0] ) );
  DFFQX2 \ImageBuffer_reg[21][2]  ( .D(n8452), .CK(clk), .Q(
        \ImageBuffer[21][2] ) );
  DFFQX2 \ImageBuffer_reg[21][0]  ( .D(n8580), .CK(clk), .Q(
        \ImageBuffer[21][0] ) );
  DFFQX2 \ImageBuffer_reg[17][2]  ( .D(n8456), .CK(clk), .Q(
        \ImageBuffer[17][2] ) );
  DFFQX2 \ImageBuffer_reg[17][0]  ( .D(n8584), .CK(clk), .Q(
        \ImageBuffer[17][0] ) );
  DFFQX2 \ImageBuffer_reg[13][2]  ( .D(n8460), .CK(clk), .Q(
        \ImageBuffer[13][2] ) );
  DFFQX2 \ImageBuffer_reg[13][0]  ( .D(n8588), .CK(clk), .Q(
        \ImageBuffer[13][0] ) );
  DFFQX2 \ImageBuffer_reg[9][2]  ( .D(n8464), .CK(clk), .Q(\ImageBuffer[9][2] ) );
  DFFQX2 \ImageBuffer_reg[9][0]  ( .D(n8592), .CK(clk), .Q(\ImageBuffer[9][0] ) );
  DFFQX2 \ImageBuffer_reg[5][2]  ( .D(n8468), .CK(clk), .Q(\ImageBuffer[5][2] ) );
  DFFQX2 \ImageBuffer_reg[5][0]  ( .D(n8596), .CK(clk), .Q(\ImageBuffer[5][0] ) );
  DFFQX2 \ImageBuffer_reg[1][2]  ( .D(n8472), .CK(clk), .Q(\ImageBuffer[1][2] ) );
  DFFQX2 \ImageBuffer_reg[1][0]  ( .D(n8600), .CK(clk), .Q(\ImageBuffer[1][0] ) );
  DFFQX2 \ImageBuffer_reg[63][2]  ( .D(n8410), .CK(clk), .Q(
        \ImageBuffer[63][2] ) );
  DFFQX2 \ImageBuffer_reg[63][0]  ( .D(n8538), .CK(clk), .Q(
        \ImageBuffer[63][0] ) );
  DFFQX2 \ImageBuffer_reg[59][2]  ( .D(n8414), .CK(clk), .Q(
        \ImageBuffer[59][2] ) );
  DFFQX2 \ImageBuffer_reg[59][0]  ( .D(n8542), .CK(clk), .Q(
        \ImageBuffer[59][0] ) );
  DFFQX2 \ImageBuffer_reg[55][0]  ( .D(n8546), .CK(clk), .Q(
        \ImageBuffer[55][0] ) );
  DFFQX2 \ImageBuffer_reg[51][2]  ( .D(n8422), .CK(clk), .Q(
        \ImageBuffer[51][2] ) );
  DFFQX2 \ImageBuffer_reg[51][0]  ( .D(n8550), .CK(clk), .Q(
        \ImageBuffer[51][0] ) );
  DFFQX2 \ImageBuffer_reg[47][0]  ( .D(n8554), .CK(clk), .Q(
        \ImageBuffer[47][0] ) );
  DFFQX2 \ImageBuffer_reg[43][0]  ( .D(n8558), .CK(clk), .Q(
        \ImageBuffer[43][0] ) );
  DFFQX2 \ImageBuffer_reg[39][2]  ( .D(n8434), .CK(clk), .Q(
        \ImageBuffer[39][2] ) );
  DFFQX2 \ImageBuffer_reg[39][0]  ( .D(n8562), .CK(clk), .Q(
        \ImageBuffer[39][0] ) );
  DFFQX2 \ImageBuffer_reg[35][0]  ( .D(n8566), .CK(clk), .Q(
        \ImageBuffer[35][0] ) );
  DFFQX2 \ImageBuffer_reg[31][0]  ( .D(n8570), .CK(clk), .Q(
        \ImageBuffer[31][0] ) );
  DFFQX2 \ImageBuffer_reg[27][2]  ( .D(n8446), .CK(clk), .Q(
        \ImageBuffer[27][2] ) );
  DFFQX2 \ImageBuffer_reg[27][0]  ( .D(n8574), .CK(clk), .Q(
        \ImageBuffer[27][0] ) );
  DFFQX2 \ImageBuffer_reg[23][2]  ( .D(n8450), .CK(clk), .Q(
        \ImageBuffer[23][2] ) );
  DFFQX2 \ImageBuffer_reg[23][0]  ( .D(n8578), .CK(clk), .Q(
        \ImageBuffer[23][0] ) );
  DFFQX2 \ImageBuffer_reg[19][2]  ( .D(n8454), .CK(clk), .Q(
        \ImageBuffer[19][2] ) );
  DFFQX2 \ImageBuffer_reg[19][0]  ( .D(n8582), .CK(clk), .Q(
        \ImageBuffer[19][0] ) );
  DFFQX2 \ImageBuffer_reg[15][2]  ( .D(n8458), .CK(clk), .Q(
        \ImageBuffer[15][2] ) );
  DFFQX2 \ImageBuffer_reg[15][0]  ( .D(n8586), .CK(clk), .Q(
        \ImageBuffer[15][0] ) );
  DFFQX2 \ImageBuffer_reg[11][2]  ( .D(n8462), .CK(clk), .Q(
        \ImageBuffer[11][2] ) );
  DFFQX2 \ImageBuffer_reg[11][0]  ( .D(n8590), .CK(clk), .Q(
        \ImageBuffer[11][0] ) );
  DFFQX2 \ImageBuffer_reg[7][2]  ( .D(n8466), .CK(clk), .Q(\ImageBuffer[7][2] ) );
  DFFQX2 \ImageBuffer_reg[7][0]  ( .D(n8594), .CK(clk), .Q(\ImageBuffer[7][0] ) );
  DFFQX2 \ImageBuffer_reg[3][2]  ( .D(n8470), .CK(clk), .Q(\ImageBuffer[3][2] ) );
  DFFQX2 \ImageBuffer_reg[3][0]  ( .D(n8598), .CK(clk), .Q(\ImageBuffer[3][0] ) );
  DFFQX2 \ImageBuffer_reg[60][2]  ( .D(n8413), .CK(clk), .Q(
        \ImageBuffer[60][2] ) );
  DFFQX2 \ImageBuffer_reg[56][0]  ( .D(n8545), .CK(clk), .Q(
        \ImageBuffer[56][0] ) );
  DFFQX2 \ImageBuffer_reg[52][2]  ( .D(n8421), .CK(clk), .Q(
        \ImageBuffer[52][2] ) );
  DFFQX2 \ImageBuffer_reg[52][0]  ( .D(n8549), .CK(clk), .Q(
        \ImageBuffer[52][0] ) );
  DFFQX2 \ImageBuffer_reg[48][2]  ( .D(n8425), .CK(clk), .Q(
        \ImageBuffer[48][2] ) );
  DFFQX2 \ImageBuffer_reg[48][0]  ( .D(n8553), .CK(clk), .Q(
        \ImageBuffer[48][0] ) );
  DFFQX2 \ImageBuffer_reg[44][0]  ( .D(n8557), .CK(clk), .Q(
        \ImageBuffer[44][0] ) );
  DFFQX2 \ImageBuffer_reg[40][0]  ( .D(n8561), .CK(clk), .Q(
        \ImageBuffer[40][0] ) );
  DFFQX2 \ImageBuffer_reg[36][2]  ( .D(n8437), .CK(clk), .Q(
        \ImageBuffer[36][2] ) );
  DFFQX2 \ImageBuffer_reg[36][0]  ( .D(n8565), .CK(clk), .Q(
        \ImageBuffer[36][0] ) );
  DFFQX2 \ImageBuffer_reg[32][0]  ( .D(n8569), .CK(clk), .Q(
        \ImageBuffer[32][0] ) );
  DFFQX2 \ImageBuffer_reg[28][0]  ( .D(n8573), .CK(clk), .Q(
        \ImageBuffer[28][0] ) );
  DFFQX2 \ImageBuffer_reg[24][2]  ( .D(n8449), .CK(clk), .Q(
        \ImageBuffer[24][2] ) );
  DFFQX2 \ImageBuffer_reg[24][0]  ( .D(n8577), .CK(clk), .Q(
        \ImageBuffer[24][0] ) );
  DFFQX2 \ImageBuffer_reg[20][2]  ( .D(n8453), .CK(clk), .Q(
        \ImageBuffer[20][2] ) );
  DFFQX2 \ImageBuffer_reg[20][0]  ( .D(n8581), .CK(clk), .Q(
        \ImageBuffer[20][0] ) );
  DFFQX2 \ImageBuffer_reg[16][2]  ( .D(n8457), .CK(clk), .Q(
        \ImageBuffer[16][2] ) );
  DFFQX2 \ImageBuffer_reg[16][0]  ( .D(n8585), .CK(clk), .Q(
        \ImageBuffer[16][0] ) );
  DFFQX2 \ImageBuffer_reg[12][2]  ( .D(n8461), .CK(clk), .Q(
        \ImageBuffer[12][2] ) );
  DFFQX2 \ImageBuffer_reg[12][0]  ( .D(n8589), .CK(clk), .Q(
        \ImageBuffer[12][0] ) );
  DFFQX2 \ImageBuffer_reg[8][2]  ( .D(n8465), .CK(clk), .Q(\ImageBuffer[8][2] ) );
  DFFQX2 \ImageBuffer_reg[8][0]  ( .D(n8593), .CK(clk), .Q(\ImageBuffer[8][0] ) );
  DFFQX2 \ImageBuffer_reg[4][2]  ( .D(n8469), .CK(clk), .Q(\ImageBuffer[4][2] ) );
  DFFQX2 \ImageBuffer_reg[4][0]  ( .D(n8597), .CK(clk), .Q(\ImageBuffer[4][0] ) );
  DFFQX2 \ImageBuffer_reg[0][2]  ( .D(n8473), .CK(clk), .Q(\ImageBuffer[0][2] ) );
  DFFQX2 \ImageBuffer_reg[0][0]  ( .D(n8601), .CK(clk), .Q(\ImageBuffer[0][0] ) );
  DFFQX2 \ImageBuffer_reg[62][2]  ( .D(n8411), .CK(clk), .Q(
        \ImageBuffer[62][2] ) );
  DFFQX2 \ImageBuffer_reg[62][0]  ( .D(n8539), .CK(clk), .Q(
        \ImageBuffer[62][0] ) );
  DFFQX2 \ImageBuffer_reg[58][2]  ( .D(n8415), .CK(clk), .Q(
        \ImageBuffer[58][2] ) );
  DFFQX2 \ImageBuffer_reg[58][0]  ( .D(n8543), .CK(clk), .Q(
        \ImageBuffer[58][0] ) );
  DFFQX2 \ImageBuffer_reg[54][2]  ( .D(n8419), .CK(clk), .Q(
        \ImageBuffer[54][2] ) );
  DFFQX2 \ImageBuffer_reg[54][0]  ( .D(n8547), .CK(clk), .Q(
        \ImageBuffer[54][0] ) );
  DFFQX2 \ImageBuffer_reg[50][0]  ( .D(n8551), .CK(clk), .Q(
        \ImageBuffer[50][0] ) );
  DFFQX2 \ImageBuffer_reg[46][0]  ( .D(n8555), .CK(clk), .Q(
        \ImageBuffer[46][0] ) );
  DFFQX2 \ImageBuffer_reg[42][0]  ( .D(n8559), .CK(clk), .Q(
        \ImageBuffer[42][0] ) );
  DFFQX2 \ImageBuffer_reg[38][2]  ( .D(n8435), .CK(clk), .Q(
        \ImageBuffer[38][2] ) );
  DFFQX2 \ImageBuffer_reg[38][0]  ( .D(n8563), .CK(clk), .Q(
        \ImageBuffer[38][0] ) );
  DFFQX2 \ImageBuffer_reg[34][0]  ( .D(n8567), .CK(clk), .Q(
        \ImageBuffer[34][0] ) );
  DFFQX2 \ImageBuffer_reg[30][0]  ( .D(n8571), .CK(clk), .Q(
        \ImageBuffer[30][0] ) );
  DFFQX2 \ImageBuffer_reg[26][2]  ( .D(n8447), .CK(clk), .Q(
        \ImageBuffer[26][2] ) );
  DFFQX2 \ImageBuffer_reg[26][0]  ( .D(n8575), .CK(clk), .Q(
        \ImageBuffer[26][0] ) );
  DFFQX2 \ImageBuffer_reg[22][2]  ( .D(n8451), .CK(clk), .Q(
        \ImageBuffer[22][2] ) );
  DFFQX2 \ImageBuffer_reg[22][0]  ( .D(n8579), .CK(clk), .Q(
        \ImageBuffer[22][0] ) );
  DFFQX2 \ImageBuffer_reg[18][2]  ( .D(n8455), .CK(clk), .Q(
        \ImageBuffer[18][2] ) );
  DFFQX2 \ImageBuffer_reg[18][0]  ( .D(n8583), .CK(clk), .Q(
        \ImageBuffer[18][0] ) );
  DFFQX2 \ImageBuffer_reg[14][2]  ( .D(n8459), .CK(clk), .Q(
        \ImageBuffer[14][2] ) );
  DFFQX2 \ImageBuffer_reg[14][0]  ( .D(n8587), .CK(clk), .Q(
        \ImageBuffer[14][0] ) );
  DFFQX2 \ImageBuffer_reg[10][2]  ( .D(n8463), .CK(clk), .Q(
        \ImageBuffer[10][2] ) );
  DFFQX2 \ImageBuffer_reg[10][0]  ( .D(n8591), .CK(clk), .Q(
        \ImageBuffer[10][0] ) );
  DFFQX2 \ImageBuffer_reg[6][2]  ( .D(n8467), .CK(clk), .Q(\ImageBuffer[6][2] ) );
  DFFQX2 \ImageBuffer_reg[6][0]  ( .D(n8595), .CK(clk), .Q(\ImageBuffer[6][0] ) );
  DFFQX2 \ImageBuffer_reg[2][2]  ( .D(n8471), .CK(clk), .Q(\ImageBuffer[2][2] ) );
  DFFQX2 \ImageBuffer_reg[2][0]  ( .D(n8599), .CK(clk), .Q(\ImageBuffer[2][0] ) );
  DFFQX2 \counter_reg[4]  ( .D(n3328), .CK(clk), .Q(N2521) );
  DFFQX1 \P0_reg[4]  ( .D(n3322), .CK(clk), .Q(N2485) );
  DFFQX1 \P0_reg[5]  ( .D(n3321), .CK(clk), .Q(N2486) );
  DFFQX1 \P0_reg[3]  ( .D(n3323), .CK(clk), .Q(N2484) );
  DFFHQX8 \P0_reg[1]  ( .D(n3325), .CK(clk), .Q(N2494) );
  DFFQX1 \IROM_A_reg[3]  ( .D(n3334), .CK(clk), .Q(n8619) );
  DFFQX1 \IROM_A_reg[4]  ( .D(n3333), .CK(clk), .Q(n8618) );
  DFFQX1 \IROM_A_reg[0]  ( .D(n3338), .CK(clk), .Q(n8622) );
  DFFQX1 \IROM_A_reg[2]  ( .D(n3335), .CK(clk), .Q(n8620) );
  DFFQX1 \IRAM_A_reg[5]  ( .D(N2522), .CK(clk), .Q(n8623) );
  DFFQX1 \IRAM_A_reg[2]  ( .D(N2519), .CK(clk), .Q(n8626) );
  DFFQX1 \IRAM_A_reg[4]  ( .D(N2521), .CK(clk), .Q(n8624) );
  EDFFX1 \IRAM_D_reg[0]  ( .D(N13071), .E(IRAM_valid), .CK(clk), .Q(n8651) );
  DFFQX1 \IROM_A_reg[1]  ( .D(n3336), .CK(clk), .Q(n8621) );
  DFFQX1 \IRAM_A_reg[0]  ( .D(n5106), .CK(clk), .Q(n8628) );
  EDFFX1 \IRAM_D_reg[1]  ( .D(N13070), .E(IRAM_valid), .CK(clk), .Q(n8650) );
  DFFQX1 \IRAM_A_reg[1]  ( .D(n5105), .CK(clk), .Q(n8627) );
  DFFQX1 \IROM_A_reg[5]  ( .D(n3337), .CK(clk), .Q(n8617) );
  DFFQX1 \IRAM_A_reg[3]  ( .D(n5104), .CK(clk), .Q(n8625) );
  EDFFX1 \IRAM_D_reg[3]  ( .D(N13068), .E(IRAM_valid), .CK(clk), .Q(n8648) );
  EDFFX1 \IRAM_D_reg[4]  ( .D(N13067), .E(IRAM_valid), .CK(clk), .Q(n8647) );
  DFFQX1 done_reg ( .D(N13653), .CK(clk), .Q(n8630) );
  EDFFX1 \IRAM_D_reg[5]  ( .D(N13066), .E(IRAM_valid), .CK(clk), .Q(n8646) );
  EDFFX1 \IRAM_D_reg[6]  ( .D(N13065), .E(IRAM_valid), .CK(clk), .Q(n8645) );
  DFFHQX8 \ImageBuffer_reg[60][0]  ( .D(n8541), .CK(clk), .Q(
        \ImageBuffer[60][0] ) );
  DFFHQX8 \ImageBuffer_reg[61][0]  ( .D(n8540), .CK(clk), .Q(
        \ImageBuffer[61][0] ) );
  DFFRX1 \state_cs_reg[0]  ( .D(state_ns[0]), .CK(clk), .RN(n8602), .Q(
        \state_cs[0] ), .QN(n8061) );
  DFFQX4 \P0_reg[2]  ( .D(n3324), .CK(clk), .Q(N2495) );
  DFFRX1 \state_cs_reg[1]  ( .D(state_ns[1]), .CK(clk), .RN(n8602), .QN(n5400)
         );
  DFFHQX4 \P0_reg[0]  ( .D(n3326), .CK(clk), .Q(N2493) );
  DFFHQX2 \ImageBuffer_reg[38][7]  ( .D(n8115), .CK(clk), .Q(
        \ImageBuffer[38][7] ) );
  DFFQX2 \ImageBuffer_reg[30][2]  ( .D(n8443), .CK(clk), .Q(
        \ImageBuffer[30][2] ) );
  DFFQX2 \ImageBuffer_reg[33][2]  ( .D(n8440), .CK(clk), .Q(
        \ImageBuffer[33][2] ) );
  DFFQX2 \ImageBuffer_reg[32][2]  ( .D(n8441), .CK(clk), .Q(
        \ImageBuffer[32][2] ) );
  DFFQX2 \ImageBuffer_reg[35][2]  ( .D(n8438), .CK(clk), .Q(
        \ImageBuffer[35][2] ) );
  DFFQX2 \ImageBuffer_reg[40][2]  ( .D(n8433), .CK(clk), .Q(
        \ImageBuffer[40][2] ) );
  DFFQX2 \ImageBuffer_reg[42][2]  ( .D(n8431), .CK(clk), .Q(
        \ImageBuffer[42][2] ) );
  DFFQX2 \ImageBuffer_reg[45][2]  ( .D(n8428), .CK(clk), .Q(
        \ImageBuffer[45][2] ) );
  DFFQX2 \ImageBuffer_reg[47][2]  ( .D(n8426), .CK(clk), .Q(
        \ImageBuffer[47][2] ) );
  DFFQX2 \ImageBuffer_reg[50][2]  ( .D(n8423), .CK(clk), .Q(
        \ImageBuffer[50][2] ) );
  DFFQX2 \ImageBuffer_reg[41][2]  ( .D(n8432), .CK(clk), .Q(
        \ImageBuffer[41][2] ) );
  DFFQX2 \ImageBuffer_reg[43][2]  ( .D(n8430), .CK(clk), .Q(
        \ImageBuffer[43][2] ) );
  DFFQX2 \ImageBuffer_reg[44][2]  ( .D(n8429), .CK(clk), .Q(
        \ImageBuffer[44][2] ) );
  DFFQX2 \ImageBuffer_reg[46][2]  ( .D(n8427), .CK(clk), .Q(
        \ImageBuffer[46][2] ) );
  DFFQX2 \ImageBuffer_reg[28][2]  ( .D(n8445), .CK(clk), .Q(
        \ImageBuffer[28][2] ) );
  DFFQX2 \ImageBuffer_reg[29][2]  ( .D(n8444), .CK(clk), .Q(
        \ImageBuffer[29][2] ) );
  DFFQX2 \ImageBuffer_reg[31][2]  ( .D(n8442), .CK(clk), .Q(
        \ImageBuffer[31][2] ) );
  DFFQX2 \ImageBuffer_reg[34][2]  ( .D(n8439), .CK(clk), .Q(
        \ImageBuffer[34][2] ) );
  DFFQX2 \ImageBuffer_reg[53][2]  ( .D(n8420), .CK(clk), .Q(
        \ImageBuffer[53][2] ) );
  DFFQX2 \ImageBuffer_reg[55][2]  ( .D(n8418), .CK(clk), .Q(
        \ImageBuffer[55][2] ) );
  DFFQX2 \ImageBuffer_reg[56][2]  ( .D(n8417), .CK(clk), .Q(
        \ImageBuffer[56][2] ) );
  AOI211X1 U3279 ( .A0(n5089), .A1(n5703), .B0(n6489), .C0(n3354), .Y(n6487)
         );
  INVX1 U3280 ( .A(n7744), .Y(n5787) );
  OAI21X1 U3281 ( .A0(n6466), .A1(n5637), .B0(n6467), .Y(n8307) );
  OAI21X1 U3282 ( .A0(n6496), .A1(n5727), .B0(n6497), .Y(n8317) );
  OAI21X1 U3283 ( .A0(n6478), .A1(n5673), .B0(n6479), .Y(n8311) );
  OAI21X1 U3284 ( .A0(n6400), .A1(n5439), .B0(n6401), .Y(n8285) );
  OAI21X1 U3285 ( .A0(n6415), .A1(n5484), .B0(n6416), .Y(n8290) );
  OAI21X1 U3286 ( .A0(n6481), .A1(n5682), .B0(n6482), .Y(n8312) );
  OAI21X1 U3287 ( .A0(n6409), .A1(n5466), .B0(n6410), .Y(n8288) );
  OAI21X1 U3288 ( .A0(n6791), .A1(n5430), .B0(n6792), .Y(n8412) );
  INVX1 U3289 ( .A(n7801), .Y(n5832) );
  OAI21X1 U3290 ( .A0(n6529), .A1(n5826), .B0(n6530), .Y(n8328) );
  AOI211XL U3291 ( .A0(n5090), .A1(n5829), .B0(n6531), .C0(n3354), .Y(n6529)
         );
  OAI21X1 U3292 ( .A0(n6777), .A1(n5979), .B0(n6778), .Y(n8409) );
  OAI21X1 U3293 ( .A0(n6642), .A1(n5574), .B0(n6643), .Y(n8364) );
  INVX1 U3294 ( .A(n7303), .Y(n5481) );
  OAI21X1 U3295 ( .A0(n6612), .A1(n5484), .B0(n6613), .Y(n8354) );
  AOI211X4 U3296 ( .A0(n5084), .A1(n5487), .B0(n6614), .C0(n3359), .Y(n6612)
         );
  OAI21X1 U3297 ( .A0(n6618), .A1(n5502), .B0(n6619), .Y(n8356) );
  AOI211X4 U3298 ( .A0(n5084), .A1(n5505), .B0(n6620), .C0(n6588), .Y(n6618)
         );
  INVX1 U3299 ( .A(n7274), .Y(n5463) );
  OAI21X1 U3300 ( .A0(n6603), .A1(n5457), .B0(n6604), .Y(n8351) );
  AOI211X4 U3301 ( .A0(n5083), .A1(n5460), .B0(n6605), .C0(n3359), .Y(n6603)
         );
  OAI21X1 U3302 ( .A0(n6672), .A1(n5664), .B0(n6673), .Y(n8374) );
  OAI21X1 U3303 ( .A0(n6678), .A1(n5682), .B0(n6679), .Y(n8376) );
  OAI21X1 U3304 ( .A0(n6690), .A1(n5718), .B0(n6691), .Y(n8380) );
  AOI211X4 U3305 ( .A0(n5084), .A1(n5721), .B0(n6692), .C0(n6588), .Y(n6690)
         );
  INVX1 U3306 ( .A(n7767), .Y(n5805) );
  OAI21X1 U3307 ( .A0(n6684), .A1(n5700), .B0(n6685), .Y(n8378) );
  AOI211X4 U3308 ( .A0(n5084), .A1(n5703), .B0(n6686), .C0(n3359), .Y(n6684)
         );
  OAI21X1 U3309 ( .A0(n6663), .A1(n5637), .B0(n6664), .Y(n8371) );
  AOI211X4 U3310 ( .A0(n5084), .A1(n5640), .B0(n6665), .C0(n6588), .Y(n6663)
         );
  OAI21X1 U3311 ( .A0(n6693), .A1(n5727), .B0(n6694), .Y(n8381) );
  AOI211X4 U3312 ( .A0(n5084), .A1(n5730), .B0(n6695), .C0(n3359), .Y(n6693)
         );
  OAI21X1 U3313 ( .A0(n6669), .A1(n5655), .B0(n6670), .Y(n8373) );
  AOI211X4 U3314 ( .A0(n5084), .A1(n5658), .B0(n6671), .C0(n6588), .Y(n6669)
         );
  OAI21X1 U3315 ( .A0(n6699), .A1(n5745), .B0(n6700), .Y(n8383) );
  AOI211X4 U3316 ( .A0(n5083), .A1(n5748), .B0(n6701), .C0(n6588), .Y(n6699)
         );
  OAI21X1 U3317 ( .A0(n6702), .A1(n5754), .B0(n6703), .Y(n8384) );
  AOI211X4 U3318 ( .A0(n5083), .A1(n5757), .B0(n6704), .C0(n3359), .Y(n6702)
         );
  INVX12 U3319 ( .A(n3497), .Y(n3498) );
  INVX4 U3320 ( .A(n3737), .Y(n3497) );
  OAI21X1 U3321 ( .A0(n6639), .A1(n5565), .B0(n6640), .Y(n8363) );
  AOI211X4 U3322 ( .A0(n5084), .A1(n5568), .B0(n6641), .C0(n3359), .Y(n6639)
         );
  OAI21X1 U3323 ( .A0(n6696), .A1(n5736), .B0(n6697), .Y(n8382) );
  AOI211X4 U3324 ( .A0(n5083), .A1(n5739), .B0(n6698), .C0(n6588), .Y(n6696)
         );
  OAI21X1 U3325 ( .A0(n6675), .A1(n5673), .B0(n6676), .Y(n8375) );
  AOI211X4 U3326 ( .A0(n5084), .A1(n5676), .B0(n6677), .C0(n3359), .Y(n6675)
         );
  OAI21X1 U3327 ( .A0(n6666), .A1(n5646), .B0(n6667), .Y(n8372) );
  AOI211X4 U3328 ( .A0(n5084), .A1(n5649), .B0(n6668), .C0(n6588), .Y(n6666)
         );
  NOR2BX1 U3329 ( .AN(n5091), .B(N2769), .Y(n5386) );
  BUFX6 U3330 ( .A(n3946), .Y(n5091) );
  OAI21X1 U3331 ( .A0(n6615), .A1(n5493), .B0(n6616), .Y(n8355) );
  AOI211X4 U3332 ( .A0(n5084), .A1(n5496), .B0(n6617), .C0(n6588), .Y(n6615)
         );
  OAI21X1 U3333 ( .A0(n6609), .A1(n5475), .B0(n6610), .Y(n8353) );
  AOI211X4 U3334 ( .A0(n5084), .A1(n5478), .B0(n6611), .C0(n3359), .Y(n6609)
         );
  OAI21X1 U3335 ( .A0(n6645), .A1(n5583), .B0(n6646), .Y(n8365) );
  AOI211X4 U3336 ( .A0(n5084), .A1(n5586), .B0(n6647), .C0(n6588), .Y(n6645)
         );
  OAI21X1 U3337 ( .A0(n6636), .A1(n5556), .B0(n6637), .Y(n8362) );
  AOI211X4 U3338 ( .A0(n5084), .A1(n5559), .B0(n6638), .C0(n3359), .Y(n6636)
         );
  OAI21X1 U3339 ( .A0(n6654), .A1(n5610), .B0(n6655), .Y(n8368) );
  AOI211X4 U3340 ( .A0(n5084), .A1(n5613), .B0(n6656), .C0(n6588), .Y(n6654)
         );
  OAI21X1 U3341 ( .A0(n6648), .A1(n5592), .B0(n6649), .Y(n8366) );
  AOI211X4 U3342 ( .A0(n5084), .A1(n5595), .B0(n6650), .C0(n3359), .Y(n6648)
         );
  OAI21X1 U3343 ( .A0(n6771), .A1(n5961), .B0(n6772), .Y(n8407) );
  AOI211X4 U3344 ( .A0(n5083), .A1(n5964), .B0(n6773), .C0(n3359), .Y(n6771)
         );
  OAI21X1 U3345 ( .A0(n6687), .A1(n5709), .B0(n6688), .Y(n8379) );
  AOI211X4 U3346 ( .A0(n5084), .A1(n5712), .B0(n6689), .C0(n6588), .Y(n6687)
         );
  OAI21X1 U3347 ( .A0(n6681), .A1(n5691), .B0(n6682), .Y(n8377) );
  AOI211X4 U3348 ( .A0(n5084), .A1(n5694), .B0(n6683), .C0(n3359), .Y(n6681)
         );
  OAI21X1 U3349 ( .A0(n6744), .A1(n5880), .B0(n6745), .Y(n8398) );
  AOI211X4 U3350 ( .A0(n5083), .A1(n5883), .B0(n6746), .C0(n6588), .Y(n6744)
         );
  OAI21X1 U3351 ( .A0(n6729), .A1(n5835), .B0(n6730), .Y(n8393) );
  AOI211X4 U3352 ( .A0(n5083), .A1(n5838), .B0(n6731), .C0(n3359), .Y(n6729)
         );
  OAI21X1 U3353 ( .A0(n6750), .A1(n5898), .B0(n6751), .Y(n8400) );
  AOI211X4 U3354 ( .A0(n5083), .A1(n5901), .B0(n6752), .C0(n6588), .Y(n6750)
         );
  OAI21X1 U3355 ( .A0(n6747), .A1(n5889), .B0(n6748), .Y(n8399) );
  AOI211X4 U3356 ( .A0(n5083), .A1(n5892), .B0(n6749), .C0(n3359), .Y(n6747)
         );
  OAI21X1 U3357 ( .A0(n6756), .A1(n5916), .B0(n6757), .Y(n8402) );
  AOI211X4 U3358 ( .A0(n5083), .A1(n5919), .B0(n6758), .C0(n6588), .Y(n6756)
         );
  OAI21X1 U3359 ( .A0(n6753), .A1(n5907), .B0(n6754), .Y(n8401) );
  AOI211X4 U3360 ( .A0(n5083), .A1(n5910), .B0(n6755), .C0(n3359), .Y(n6753)
         );
  OAI21X1 U3361 ( .A0(n6711), .A1(n5781), .B0(n6712), .Y(n8387) );
  AOI211X4 U3362 ( .A0(n5083), .A1(n5784), .B0(n6713), .C0(n6588), .Y(n6711)
         );
  OAI21X1 U3363 ( .A0(n6630), .A1(n5538), .B0(n6631), .Y(n8360) );
  AOI211X4 U3364 ( .A0(n5084), .A1(n5541), .B0(n6632), .C0(n3359), .Y(n6630)
         );
  OAI21X1 U3365 ( .A0(n6720), .A1(n5808), .B0(n6721), .Y(n8390) );
  AOI211X4 U3366 ( .A0(n5083), .A1(n5811), .B0(n6722), .C0(n6588), .Y(n6720)
         );
  OAI21X1 U3367 ( .A0(n6621), .A1(n5511), .B0(n6622), .Y(n8357) );
  AOI211X4 U3368 ( .A0(n5084), .A1(n5514), .B0(n6623), .C0(n3359), .Y(n6621)
         );
  OAI21X1 U3369 ( .A0(n6726), .A1(n5826), .B0(n6727), .Y(n8392) );
  AOI211X4 U3370 ( .A0(n5083), .A1(n5829), .B0(n6728), .C0(n6588), .Y(n6726)
         );
  OAI21X1 U3371 ( .A0(n6708), .A1(n5772), .B0(n6709), .Y(n8386) );
  AOI211X4 U3372 ( .A0(n5083), .A1(n5775), .B0(n6710), .C0(n3359), .Y(n6708)
         );
  OAI21X1 U3373 ( .A0(n6732), .A1(n5844), .B0(n6733), .Y(n8394) );
  AOI211X4 U3374 ( .A0(n5083), .A1(n5847), .B0(n6734), .C0(n6588), .Y(n6732)
         );
  OAI21X1 U3375 ( .A0(n6714), .A1(n5790), .B0(n6715), .Y(n8388) );
  AOI211X4 U3376 ( .A0(n5083), .A1(n5793), .B0(n6716), .C0(n3359), .Y(n6714)
         );
  OAI21X1 U3377 ( .A0(n6738), .A1(n5862), .B0(n6739), .Y(n8396) );
  AOI211X4 U3378 ( .A0(n5083), .A1(n5865), .B0(n6740), .C0(n6588), .Y(n6738)
         );
  OAI21X1 U3379 ( .A0(n6723), .A1(n5817), .B0(n6724), .Y(n8391) );
  AOI211X4 U3380 ( .A0(n5083), .A1(n5820), .B0(n6725), .C0(n3359), .Y(n6723)
         );
  OAI21X1 U3381 ( .A0(n6660), .A1(n5628), .B0(n6661), .Y(n8370) );
  AOI211X4 U3382 ( .A0(n5084), .A1(n5631), .B0(n6662), .C0(n6588), .Y(n6660)
         );
  OAI21X1 U3383 ( .A0(n6735), .A1(n5853), .B0(n6736), .Y(n8395) );
  AOI211X4 U3384 ( .A0(n5083), .A1(n5856), .B0(n6737), .C0(n3359), .Y(n6735)
         );
  OAI21X1 U3385 ( .A0(n6633), .A1(n5547), .B0(n6634), .Y(n8361) );
  AOI211X4 U3386 ( .A0(n5084), .A1(n5550), .B0(n6635), .C0(n6588), .Y(n6633)
         );
  OAI21X1 U3387 ( .A0(n6624), .A1(n5520), .B0(n6625), .Y(n8358) );
  AOI211X4 U3388 ( .A0(n5084), .A1(n5523), .B0(n6626), .C0(n3359), .Y(n6624)
         );
  OAI21X1 U3389 ( .A0(n6705), .A1(n5763), .B0(n6706), .Y(n8385) );
  AOI211X4 U3390 ( .A0(n5083), .A1(n5766), .B0(n6707), .C0(n6588), .Y(n6705)
         );
  BUFX4 U3391 ( .A(n3942), .Y(n3936) );
  OAI21X1 U3392 ( .A0(n6600), .A1(n5448), .B0(n6601), .Y(n8350) );
  AOI211X4 U3393 ( .A0(n5084), .A1(n5451), .B0(n6602), .C0(n3359), .Y(n6600)
         );
  OAI21X1 U3394 ( .A0(n6762), .A1(n5934), .B0(n6763), .Y(n8404) );
  AOI211X4 U3395 ( .A0(n5083), .A1(n5937), .B0(n6764), .C0(n6588), .Y(n6762)
         );
  OAI21X1 U3396 ( .A0(n6759), .A1(n5925), .B0(n6760), .Y(n8403) );
  AOI211X4 U3397 ( .A0(n5083), .A1(n5928), .B0(n6761), .C0(n3359), .Y(n6759)
         );
  OAI21X1 U3398 ( .A0(n6768), .A1(n5952), .B0(n6769), .Y(n8406) );
  AOI211X4 U3399 ( .A0(n5083), .A1(n5955), .B0(n6770), .C0(n6588), .Y(n6768)
         );
  OAI21X1 U3400 ( .A0(n6765), .A1(n5943), .B0(n6766), .Y(n8405) );
  AOI211X4 U3401 ( .A0(n5083), .A1(n5946), .B0(n6767), .C0(n3359), .Y(n6765)
         );
  OAI21X1 U3402 ( .A0(n6606), .A1(n5466), .B0(n6607), .Y(n8352) );
  AOI211X4 U3403 ( .A0(n5084), .A1(n5469), .B0(n6608), .C0(n6588), .Y(n6606)
         );
  OAI21X1 U3404 ( .A0(n6774), .A1(n5970), .B0(n6775), .Y(n8408) );
  AOI211X4 U3405 ( .A0(n5083), .A1(n5973), .B0(n6776), .C0(n3359), .Y(n6774)
         );
  OAI21X1 U3406 ( .A0(n6627), .A1(n5529), .B0(n6628), .Y(n8359) );
  AOI211X4 U3407 ( .A0(n5084), .A1(n5532), .B0(n6629), .C0(n6588), .Y(n6627)
         );
  OAI21X1 U3408 ( .A0(n6651), .A1(n5601), .B0(n6652), .Y(n8367) );
  AOI211X4 U3409 ( .A0(n5084), .A1(n5604), .B0(n6653), .C0(n6588), .Y(n6651)
         );
  OAI21X1 U3410 ( .A0(n6657), .A1(n5619), .B0(n6658), .Y(n8369) );
  AOI211X4 U3411 ( .A0(n5084), .A1(n5622), .B0(n6659), .C0(n3359), .Y(n6657)
         );
  INVX1 U3412 ( .A(n7655), .Y(n5724) );
  INVX1 U3413 ( .A(n7325), .Y(n5490) );
  OAI222X4 U3414 ( .A0(n5534), .A1(n5017), .B0(n5535), .B1(n6787), .C0(n5536), 
        .C1(n5024), .Y(n6826) );
  INVX1 U3415 ( .A(n7386), .Y(n5535) );
  OAI222XL U3416 ( .A0(n5750), .A1(n6983), .B0(n5751), .B1(n5034), .C0(n5752), 
        .C1(n6985), .Y(n7096) );
  INVX3 U3417 ( .A(n7691), .Y(n5750) );
  INVX1 U3418 ( .A(n7628), .Y(n5706) );
  INVX1 U3419 ( .A(n7452), .Y(n5580) );
  INVX1 U3420 ( .A(n7425), .Y(n5562) );
  INVX3 U3421 ( .A(n7732), .Y(n5777) );
  INVX3 U3422 ( .A(n7758), .Y(n5795) );
  OAI222X4 U3423 ( .A0(n5786), .A1(n4990), .B0(n5787), .B1(n4992), .C0(n5788), 
        .C1(n4996), .Y(n6516) );
  INVX3 U3424 ( .A(n7745), .Y(n5786) );
  OAI222X4 U3425 ( .A0(n5606), .A1(n5016), .B0(n5607), .B1(n5020), .C0(n5608), 
        .C1(n5023), .Y(n6850) );
  INVX1 U3426 ( .A(n7486), .Y(n5607) );
  INVX3 U3427 ( .A(n7557), .Y(n5651) );
  ADDHX4 U3428 ( .A(n5127), .B(\r2549/carry[3] ), .CO(\r2549/carry[4] ), .S(
        N2490) );
  ADDHX4 U3429 ( .A(N2495), .B(\r2549/carry[2] ), .CO(\r2549/carry[3] ), .S(
        N2489) );
  INVX3 U3430 ( .A(n7891), .Y(n5894) );
  OAI222X4 U3431 ( .A0(n5831), .A1(n4979), .B0(n5832), .B1(n4980), .C0(n5833), 
        .C1(n4984), .Y(n6333) );
  INVX3 U3432 ( .A(n7802), .Y(n5831) );
  INVX3 U3433 ( .A(n7792), .Y(n5822) );
  CLKBUFX8 U3434 ( .A(N2501), .Y(n3487) );
  AOI211XL U3435 ( .A0(n5089), .A1(n5983), .B0(n6582), .C0(n3356), .Y(n6580)
         );
  AOI211XL U3436 ( .A0(n5089), .A1(n5568), .B0(n6444), .C0(n3356), .Y(n6442)
         );
  AOI211XL U3437 ( .A0(n5089), .A1(n5730), .B0(n6498), .C0(n3354), .Y(n6496)
         );
  AOI211XL U3438 ( .A0(n5089), .A1(n5712), .B0(n6492), .C0(n3355), .Y(n6490)
         );
  AOI211XL U3439 ( .A0(n5089), .A1(n5694), .B0(n6486), .C0(n3356), .Y(n6484)
         );
  AOI211XL U3440 ( .A0(n5089), .A1(n5676), .B0(n6480), .C0(n3354), .Y(n6478)
         );
  AOI211XL U3441 ( .A0(n5089), .A1(n5667), .B0(n6477), .C0(n3355), .Y(n6475)
         );
  AOI211XL U3442 ( .A0(n5089), .A1(n5640), .B0(n6468), .C0(n3354), .Y(n6466)
         );
  AOI211XL U3443 ( .A0(n5089), .A1(n5622), .B0(n6462), .C0(n3355), .Y(n6460)
         );
  AOI211XL U3444 ( .A0(n5089), .A1(n5523), .B0(n6429), .C0(n3356), .Y(n6427)
         );
  AOI211XL U3445 ( .A0(n5089), .A1(n5550), .B0(n6438), .C0(n3356), .Y(n6436)
         );
  AOI211XL U3446 ( .A0(n5089), .A1(n5514), .B0(n6426), .C0(n3355), .Y(n6424)
         );
  AOI211XL U3447 ( .A0(n5089), .A1(n5721), .B0(n6495), .C0(n3356), .Y(n6493)
         );
  AOI211XL U3448 ( .A0(n5089), .A1(n5685), .B0(n6483), .C0(n3354), .Y(n6481)
         );
  AOI211XL U3449 ( .A0(n5089), .A1(n5541), .B0(n6435), .C0(n3355), .Y(n6433)
         );
  AOI211XL U3450 ( .A0(n5089), .A1(n5487), .B0(n6417), .C0(n3354), .Y(n6415)
         );
  BUFX8 U3451 ( .A(n5089), .Y(n5090) );
  AND2X2 U3452 ( .A(n5161), .B(n5171), .Y(n5168) );
  OAI222X4 U3453 ( .A0(n5723), .A1(n5015), .B0(n5724), .B1(n5018), .C0(n5725), 
        .C1(n5023), .Y(n6889) );
  INVX3 U3454 ( .A(n7657), .Y(n5723) );
  BUFX12 U3455 ( .A(n3546), .Y(n5114) );
  XNOR2X2 U3456 ( .A(n3747), .B(n5118), .Y(n3546) );
  OAI31X2 U3457 ( .A0(n5185), .A1(n5184), .A2(n5183), .B0(n5182), .Y(N2696) );
  AOI211X2 U3458 ( .A0(n5181), .A1(n5180), .B0(n5179), .C0(n5178), .Y(n5183)
         );
  INVX3 U3459 ( .A(n7531), .Y(n5633) );
  CLKBUFX3 U3460 ( .A(n3928), .Y(n3339) );
  BUFX4 U3461 ( .A(n3928), .Y(n3340) );
  BUFX4 U3462 ( .A(n3928), .Y(n3341) );
  BUFX12 U3463 ( .A(N2780), .Y(n4866) );
  INVX2 U3464 ( .A(n4866), .Y(n6985) );
  CLKINVX1 U3465 ( .A(n4866), .Y(n5155) );
  AO21X4 U3466 ( .A0(n6985), .A1(n5324), .B0(n5077), .Y(n5159) );
  OAI222X4 U3467 ( .A0(n5435), .A1(n4978), .B0(n5436), .B1(n4982), .C0(n5437), 
        .C1(n4983), .Y(n6201) );
  INVX3 U3468 ( .A(n7233), .Y(n5435) );
  AO21X4 U3469 ( .A0(n6985), .A1(n3345), .B0(N2772), .Y(n5190) );
  OAI211X2 U3470 ( .A0(n3345), .A1(n6985), .B0(n5190), .C0(n5200), .Y(n5192)
         );
  OAI222X4 U3471 ( .A0(n5462), .A1(n6391), .B0(n5463), .B1(n4993), .C0(n5464), 
        .C1(n4995), .Y(n6408) );
  INVX3 U3472 ( .A(n7276), .Y(n5462) );
  INVX3 U3473 ( .A(n7262), .Y(n5453) );
  INVX3 U3474 ( .A(n7289), .Y(n5471) );
  INVX3 U3475 ( .A(n7247), .Y(n5444) );
  INVX3 U3476 ( .A(n7217), .Y(n5426) );
  BUFX20 U3477 ( .A(n5116), .Y(n3747) );
  CLKINVX4 U3478 ( .A(n5377), .Y(n5398) );
  NOR3BX1 U3479 ( .AN(n5392), .B(n5391), .C(n5376), .Y(n5377) );
  BUFX20 U3480 ( .A(n3508), .Y(n3342) );
  CLKBUFX20 U3481 ( .A(n3508), .Y(n3343) );
  CLKINVX8 U3482 ( .A(n3505), .Y(n3508) );
  INVX3 U3483 ( .A(n8026), .Y(n5990) );
  OAI222X4 U3484 ( .A0(n5507), .A1(n5017), .B0(n5508), .B1(n6787), .C0(n5509), 
        .C1(n5024), .Y(n6817) );
  INVX3 U3485 ( .A(n7354), .Y(n5507) );
  OAI222X4 U3486 ( .A0(n5489), .A1(n5017), .B0(n5490), .B1(n6787), .C0(n5491), 
        .C1(n5024), .Y(n6811) );
  INVX3 U3487 ( .A(n7328), .Y(n5489) );
  OAI222X4 U3488 ( .A0(n5480), .A1(n5017), .B0(n5481), .B1(n6787), .C0(n5482), 
        .C1(n5024), .Y(n6808) );
  INVX3 U3489 ( .A(n7306), .Y(n5480) );
  BUFX12 U3490 ( .A(n7181), .Y(n3344) );
  BUFX6 U3491 ( .A(n5191), .Y(n3345) );
  OAI21X4 U3492 ( .A0(n6741), .A1(n5871), .B0(n6742), .Y(n8397) );
  NAND2X4 U3493 ( .A(n5041), .B(n4930), .Y(n5871) );
  AOI211X4 U3494 ( .A0(n5083), .A1(n5874), .B0(n6743), .C0(n3359), .Y(n6741)
         );
  OAI21X1 U3495 ( .A0(n6717), .A1(n5799), .B0(n6718), .Y(n8389) );
  AOI211X4 U3496 ( .A0(n5083), .A1(n5802), .B0(n6719), .C0(n6588), .Y(n6717)
         );
  BUFX8 U3497 ( .A(n3507), .Y(n3346) );
  CLKBUFX20 U3498 ( .A(n3507), .Y(n3347) );
  INVX4 U3499 ( .A(n3505), .Y(n3507) );
  OAI21X4 U3500 ( .A0(n6594), .A1(n5430), .B0(n6595), .Y(n8348) );
  AOI211X4 U3501 ( .A0(n5084), .A1(n5433), .B0(n6596), .C0(n3359), .Y(n6594)
         );
  OAI21X4 U3502 ( .A0(n6597), .A1(n5439), .B0(n6598), .Y(n8349) );
  AOI211X4 U3503 ( .A0(n5084), .A1(n5442), .B0(n6599), .C0(n6588), .Y(n6597)
         );
  OAI21X4 U3504 ( .A0(n6591), .A1(n5421), .B0(n6592), .Y(n8347) );
  AOI211X4 U3505 ( .A0(n5084), .A1(n5424), .B0(n6593), .C0(n6588), .Y(n6591)
         );
  OAI21X1 U3506 ( .A0(n6584), .A1(n5408), .B0(n6585), .Y(n8346) );
  AOI211X4 U3507 ( .A0(n5084), .A1(n5412), .B0(n6587), .C0(n3359), .Y(n6584)
         );
  BUFX12 U3508 ( .A(n4124), .Y(n4125) );
  BUFX12 U3509 ( .A(n8062), .Y(n3348) );
  BUFX6 U3510 ( .A(n3937), .Y(n3935) );
  CLKBUFX4 U3511 ( .A(n3942), .Y(n3937) );
  INVX3 U3512 ( .A(n7768), .Y(n5804) );
  OAI32X4 U3513 ( .A0(n7762), .A1(n5057), .A2(n7763), .B0(n3352), .B1(n7769), 
        .Y(n7768) );
  INVX2 U3514 ( .A(n4871), .Y(n5277) );
  CLKINVX1 U3515 ( .A(n4871), .Y(n5309) );
  CLKINVX2 U3516 ( .A(n4871), .Y(n6589) );
  CLKBUFX4 U3517 ( .A(n6589), .Y(n5003) );
  MX4X2 U3518 ( .A(n3839), .B(n3829), .C(n3834), .D(n3824), .S0(N2492), .S1(
        N2491), .Y(N2762) );
  BUFX12 U3519 ( .A(N2762), .Y(n4871) );
  NOR2X2 U3520 ( .A(n5187), .B(n5096), .Y(n5184) );
  INVX3 U3521 ( .A(n7857), .Y(n5867) );
  OAI32X4 U3522 ( .A0(n7849), .A1(n5058), .A2(n7850), .B0(n3351), .B1(n7856), 
        .Y(n7857) );
  INVX3 U3523 ( .A(n7831), .Y(n5849) );
  OAI32X4 U3524 ( .A0(n7822), .A1(n5058), .A2(n7823), .B0(n3352), .B1(n7830), 
        .Y(n7831) );
  MX4X2 U3525 ( .A(\ImageBuffer[24][0] ), .B(\ImageBuffer[25][0] ), .C(
        \ImageBuffer[26][0] ), .D(\ImageBuffer[27][0] ), .S0(n4114), .S1(n4130), .Y(n3959) );
  MX4XL U3526 ( .A(\ImageBuffer[40][0] ), .B(\ImageBuffer[41][0] ), .C(
        \ImageBuffer[42][0] ), .D(\ImageBuffer[43][0] ), .S0(n4114), .S1(n3753), .Y(n3955) );
  MX4XL U3527 ( .A(\ImageBuffer[32][0] ), .B(\ImageBuffer[33][0] ), .C(
        \ImageBuffer[34][0] ), .D(\ImageBuffer[35][0] ), .S0(n4114), .S1(n4134), .Y(n3957) );
  BUFX20 U3528 ( .A(n4113), .Y(n4114) );
  INVX12 U3529 ( .A(n3469), .Y(n3349) );
  INVX12 U3530 ( .A(n3469), .Y(n3350) );
  BUFX12 U3531 ( .A(n6385), .Y(n3469) );
  INVX3 U3532 ( .A(n7933), .Y(n5921) );
  OAI32X4 U3533 ( .A0(n7920), .A1(n5058), .A2(n7921), .B0(n3352), .B1(n7932), 
        .Y(n7933) );
  BUFX12 U3534 ( .A(n3365), .Y(n3351) );
  BUFX12 U3535 ( .A(n3365), .Y(n3352) );
  AND2XL U3536 ( .A(n8030), .B(n8028), .Y(n3365) );
  CLKBUFX20 U3537 ( .A(n3937), .Y(n3939) );
  AOI31X2 U3538 ( .A0(n5177), .A1(n5176), .A2(n5175), .B0(n5174), .Y(n5181) );
  INVX20 U3539 ( .A(n7304), .Y(n7192) );
  CLKBUFX2 U3540 ( .A(n7192), .Y(n5051) );
  NAND2X4 U3541 ( .A(n8028), .B(n8029), .Y(n7304) );
  INVX3 U3542 ( .A(n7973), .Y(n5948) );
  OAI32X4 U3543 ( .A0(n7965), .A1(n5058), .A2(n7966), .B0(n3351), .B1(n7974), 
        .Y(n7973) );
  INVX3 U3544 ( .A(n7985), .Y(n5957) );
  OAI32X4 U3545 ( .A0(n7978), .A1(n5058), .A2(n7979), .B0(n3351), .B1(n7986), 
        .Y(n7985) );
  CLKBUFX8 U3546 ( .A(n4299), .Y(n4297) );
  INVX3 U3547 ( .A(n8008), .Y(n5975) );
  OAI32X4 U3548 ( .A0(n8002), .A1(n5058), .A2(n8003), .B0(n3352), .B1(n8009), 
        .Y(n8008) );
  OAI221X1 U3549 ( .A0(n5117), .A1(n3348), .B0(n3490), .B1(n8063), .C0(n8070), 
        .Y(N2512) );
  NAND2BX2 U3550 ( .AN(n8074), .B(n8073), .Y(n8062) );
  MX4X2 U3551 ( .A(n4478), .B(n4468), .C(n4473), .D(n4463), .S0(N2510), .S1(
        N2509), .Y(N2742) );
  MX4X1 U3552 ( .A(n4477), .B(n4475), .C(n4476), .D(n4474), .S0(n3503), .S1(
        n3495), .Y(n4478) );
  MX4X4 U3553 ( .A(n4196), .B(n4186), .C(n4191), .D(n4181), .S0(N2504), .S1(
        N2503), .Y(N2771) );
  CLKINVX20 U3554 ( .A(n6390), .Y(n3353) );
  CLKINVX20 U3555 ( .A(n3353), .Y(n3354) );
  CLKINVX20 U3556 ( .A(n3353), .Y(n3355) );
  CLKINVX20 U3557 ( .A(n3353), .Y(n3356) );
  INVX12 U3558 ( .A(n8020), .Y(n3357) );
  INVX12 U3559 ( .A(n8020), .Y(n3358) );
  AND3X8 U3560 ( .A(n3440), .B(n3441), .C(n3442), .Y(n8020) );
  AND3X8 U3561 ( .A(n3566), .B(n3567), .C(n3568), .Y(n6187) );
  NAND2X2 U3562 ( .A(N2743), .B(n4943), .Y(n3566) );
  NAND2X2 U3563 ( .A(N2751), .B(n5988), .Y(n3568) );
  BUFX16 U3564 ( .A(n4111), .Y(n4118) );
  BUFX20 U3565 ( .A(n4111), .Y(n4119) );
  CLKBUFX4 U3566 ( .A(n5116), .Y(n3748) );
  CLKINVX20 U3567 ( .A(n5117), .Y(n5116) );
  OAI211XL U3568 ( .A0(n5324), .A1(n6985), .B0(n5159), .C0(n5168), .Y(n5160)
         );
  INVX4 U3569 ( .A(N2507), .Y(n3494) );
  OAI221X4 U3570 ( .A0(n5115), .A1(n8076), .B0(n5112), .B1(n8077), .C0(n8083), 
        .Y(N2507) );
  CLKBUFX4 U3571 ( .A(n4120), .Y(n4111) );
  MX4XL U3572 ( .A(\ImageBuffer[20][3] ), .B(\ImageBuffer[21][3] ), .C(
        \ImageBuffer[22][3] ), .D(\ImageBuffer[23][3] ), .S0(n4116), .S1(n3748), .Y(n4020) );
  MX4X4 U3573 ( .A(\ImageBuffer[16][3] ), .B(\ImageBuffer[17][3] ), .C(
        \ImageBuffer[18][3] ), .D(\ImageBuffer[19][3] ), .S0(n4116), .S1(n4132), .Y(n4021) );
  BUFX20 U3574 ( .A(n4112), .Y(n4116) );
  BUFX20 U3575 ( .A(n3922), .Y(n3929) );
  BUFX8 U3576 ( .A(n3932), .Y(n3922) );
  INVX16 U3577 ( .A(n6780), .Y(n3359) );
  AND3X8 U3578 ( .A(n3444), .B(n3445), .C(n3446), .Y(n6780) );
  CLKBUFX8 U3579 ( .A(n3947), .Y(n3360) );
  CLKBUFX8 U3580 ( .A(n3947), .Y(n3361) );
  MX4X2 U3581 ( .A(n4067), .B(n4057), .C(n4062), .D(n4052), .S0(N2498), .S1(
        N2497), .Y(n3947) );
  BUFX8 U3582 ( .A(N2508), .Y(n3362) );
  OAI221X4 U3583 ( .A0(n5127), .A1(n8076), .B0(n5109), .B1(n8077), .C0(n8082), 
        .Y(N2508) );
  CLKINVX12 U3584 ( .A(n3504), .Y(n3472) );
  OAI31X2 U3585 ( .A0(n5275), .A1(n5274), .A2(n5273), .B0(n5272), .Y(N2702) );
  AOI211X2 U3586 ( .A0(n5271), .A1(n5270), .B0(n5269), .C0(n5268), .Y(n5273)
         );
  CLKINVX20 U3587 ( .A(n5109), .Y(n5108) );
  NOR2BX4 U3588 ( .AN(N2781), .B(N2765), .Y(n5222) );
  CLKINVX12 U3589 ( .A(n3572), .Y(N2765) );
  OAI21X4 U3590 ( .A0(n6025), .A1(n5502), .B0(n6026), .Y(n8164) );
  AOI211X4 U3591 ( .A0(n5095), .A1(n5505), .B0(n6027), .C0(n5996), .Y(n6025)
         );
  OAI21X4 U3592 ( .A0(n6010), .A1(n5457), .B0(n6011), .Y(n8159) );
  AOI211X4 U3593 ( .A0(n5096), .A1(n5460), .B0(n6012), .C0(n3364), .Y(n6010)
         );
  OAI21X4 U3594 ( .A0(n6076), .A1(n5655), .B0(n6077), .Y(n8181) );
  AOI211X4 U3595 ( .A0(n5095), .A1(n5658), .B0(n6078), .C0(n5996), .Y(n6076)
         );
  OAI21X4 U3596 ( .A0(n6046), .A1(n5565), .B0(n6047), .Y(n8171) );
  AOI211X4 U3597 ( .A0(n5095), .A1(n5568), .B0(n6048), .C0(n3364), .Y(n6046)
         );
  OAI21X4 U3598 ( .A0(n6016), .A1(n5475), .B0(n6017), .Y(n8161) );
  AOI211X4 U3599 ( .A0(n5095), .A1(n5478), .B0(n6018), .C0(n5996), .Y(n6016)
         );
  OAI21X4 U3600 ( .A0(n6151), .A1(n5880), .B0(n6152), .Y(n8206) );
  AOI211X4 U3601 ( .A0(n5094), .A1(n5883), .B0(n6153), .C0(n3364), .Y(n6151)
         );
  OAI21X4 U3602 ( .A0(n6160), .A1(n5907), .B0(n6161), .Y(n8209) );
  AOI211X4 U3603 ( .A0(n5094), .A1(n5910), .B0(n6162), .C0(n5996), .Y(n6160)
         );
  OAI21X4 U3604 ( .A0(n6157), .A1(n5898), .B0(n6158), .Y(n8208) );
  AOI211X4 U3605 ( .A0(n5094), .A1(n5901), .B0(n6159), .C0(n3364), .Y(n6157)
         );
  OAI21X4 U3606 ( .A0(n6001), .A1(n5430), .B0(n6002), .Y(n8156) );
  AOI211X4 U3607 ( .A0(n5096), .A1(n5433), .B0(n6003), .C0(n5996), .Y(n6001)
         );
  OAI21X4 U3608 ( .A0(n6178), .A1(n5961), .B0(n6179), .Y(n8215) );
  AOI211X4 U3609 ( .A0(n5094), .A1(n5964), .B0(n6180), .C0(n3364), .Y(n6178)
         );
  OAI21X4 U3610 ( .A0(n6052), .A1(n5583), .B0(n6053), .Y(n8173) );
  AOI211X4 U3611 ( .A0(n5095), .A1(n5586), .B0(n6054), .C0(n5996), .Y(n6052)
         );
  OAI21X4 U3612 ( .A0(n6061), .A1(n5610), .B0(n6062), .Y(n8176) );
  AOI211X4 U3613 ( .A0(n5095), .A1(n5613), .B0(n6063), .C0(n3364), .Y(n6061)
         );
  OAI21X4 U3614 ( .A0(n6154), .A1(n5889), .B0(n6155), .Y(n8207) );
  AOI211X4 U3615 ( .A0(n5094), .A1(n5892), .B0(n6156), .C0(n5996), .Y(n6154)
         );
  OAI21X4 U3616 ( .A0(n6127), .A1(n5808), .B0(n6128), .Y(n8198) );
  AOI211X4 U3617 ( .A0(n5094), .A1(n5811), .B0(n6129), .C0(n3364), .Y(n6127)
         );
  OAI21X4 U3618 ( .A0(n6163), .A1(n5916), .B0(n6164), .Y(n8210) );
  AOI211X4 U3619 ( .A0(n5094), .A1(n5919), .B0(n6165), .C0(n5996), .Y(n6163)
         );
  OAI21X4 U3620 ( .A0(n6034), .A1(n5529), .B0(n6035), .Y(n8167) );
  AOI211X4 U3621 ( .A0(n5095), .A1(n5532), .B0(n6036), .C0(n3364), .Y(n6034)
         );
  OAI21X4 U3622 ( .A0(n6136), .A1(n5835), .B0(n6137), .Y(n8201) );
  AOI211X4 U3623 ( .A0(n5094), .A1(n5838), .B0(n6138), .C0(n5996), .Y(n6136)
         );
  OAI21X4 U3624 ( .A0(n6166), .A1(n5925), .B0(n6167), .Y(n8211) );
  AOI211X4 U3625 ( .A0(n5094), .A1(n5928), .B0(n6168), .C0(n3364), .Y(n6166)
         );
  BUFX6 U3626 ( .A(N2512), .Y(n3363) );
  OAI21X4 U3627 ( .A0(n6169), .A1(n5934), .B0(n6170), .Y(n8212) );
  AOI211X4 U3628 ( .A0(n5094), .A1(n5937), .B0(n6171), .C0(n5996), .Y(n6169)
         );
  OAI21X4 U3629 ( .A0(n6172), .A1(n5943), .B0(n6173), .Y(n8213) );
  AOI211X4 U3630 ( .A0(n5094), .A1(n5946), .B0(n6174), .C0(n3364), .Y(n6172)
         );
  OAI21X4 U3631 ( .A0(n6175), .A1(n5952), .B0(n6176), .Y(n8214) );
  AOI211X4 U3632 ( .A0(n5094), .A1(n5955), .B0(n6177), .C0(n5996), .Y(n6175)
         );
  OAI21X4 U3633 ( .A0(n6181), .A1(n5970), .B0(n6182), .Y(n8216) );
  AOI211X4 U3634 ( .A0(n5094), .A1(n5973), .B0(n6183), .C0(n3364), .Y(n6181)
         );
  OAI21X4 U3635 ( .A0(n6022), .A1(n5493), .B0(n6023), .Y(n8163) );
  AOI211X4 U3636 ( .A0(n5095), .A1(n5496), .B0(n6024), .C0(n5996), .Y(n6022)
         );
  OAI21X4 U3637 ( .A0(n6040), .A1(n5547), .B0(n6041), .Y(n8169) );
  AOI211X4 U3638 ( .A0(n5095), .A1(n5550), .B0(n6042), .C0(n3364), .Y(n6040)
         );
  OAI21X4 U3639 ( .A0(n6031), .A1(n5520), .B0(n6032), .Y(n8166) );
  AOI211X4 U3640 ( .A0(n5095), .A1(n5523), .B0(n6033), .C0(n5996), .Y(n6031)
         );
  OAI21X4 U3641 ( .A0(n6094), .A1(n5709), .B0(n6095), .Y(n8187) );
  AOI211X4 U3642 ( .A0(n5095), .A1(n5712), .B0(n6096), .C0(n3364), .Y(n6094)
         );
  OAI21X4 U3643 ( .A0(n6088), .A1(n5691), .B0(n6089), .Y(n8185) );
  AOI211X4 U3644 ( .A0(n5095), .A1(n5694), .B0(n6090), .C0(n5996), .Y(n6088)
         );
  OAI21X4 U3645 ( .A0(n6091), .A1(n5700), .B0(n6092), .Y(n8186) );
  AOI211X4 U3646 ( .A0(n5095), .A1(n5703), .B0(n6093), .C0(n3364), .Y(n6091)
         );
  OAI21X4 U3647 ( .A0(n6055), .A1(n5592), .B0(n6056), .Y(n8174) );
  AOI211X4 U3648 ( .A0(n5095), .A1(n5595), .B0(n6057), .C0(n5996), .Y(n6055)
         );
  OAI21X4 U3649 ( .A0(n6100), .A1(n5727), .B0(n6101), .Y(n8189) );
  AOI211X4 U3650 ( .A0(n5095), .A1(n5730), .B0(n6102), .C0(n3364), .Y(n6100)
         );
  OAI21X4 U3651 ( .A0(n6064), .A1(n5619), .B0(n6065), .Y(n8177) );
  AOI211X4 U3652 ( .A0(n5095), .A1(n5622), .B0(n6066), .C0(n5996), .Y(n6064)
         );
  OAI21X4 U3653 ( .A0(n6058), .A1(n5601), .B0(n6059), .Y(n8175) );
  AOI211X4 U3654 ( .A0(n5095), .A1(n5604), .B0(n6060), .C0(n3364), .Y(n6058)
         );
  OAI21X4 U3655 ( .A0(n6019), .A1(n5484), .B0(n6020), .Y(n8162) );
  AOI211X4 U3656 ( .A0(n5095), .A1(n5487), .B0(n6021), .C0(n5996), .Y(n6019)
         );
  OAI21X4 U3657 ( .A0(n6049), .A1(n5574), .B0(n6050), .Y(n8172) );
  AOI211X4 U3658 ( .A0(n5095), .A1(n5577), .B0(n6051), .C0(n3364), .Y(n6049)
         );
  OAI21X4 U3659 ( .A0(n6037), .A1(n5538), .B0(n6038), .Y(n8168) );
  AOI211X4 U3660 ( .A0(n5095), .A1(n5541), .B0(n6039), .C0(n5996), .Y(n6037)
         );
  OAI21X4 U3661 ( .A0(n6070), .A1(n5637), .B0(n6071), .Y(n8179) );
  AOI211X4 U3662 ( .A0(n5095), .A1(n5640), .B0(n6072), .C0(n3364), .Y(n6070)
         );
  OAI21X4 U3663 ( .A0(n6085), .A1(n5682), .B0(n6086), .Y(n8184) );
  AOI211X4 U3664 ( .A0(n5095), .A1(n5685), .B0(n6087), .C0(n5996), .Y(n6085)
         );
  OAI21X4 U3665 ( .A0(n6028), .A1(n5511), .B0(n6029), .Y(n8165) );
  AOI211X4 U3666 ( .A0(n5095), .A1(n5514), .B0(n6030), .C0(n3364), .Y(n6028)
         );
  OAI21X4 U3667 ( .A0(n6109), .A1(n5754), .B0(n6110), .Y(n8192) );
  AOI211X4 U3668 ( .A0(n5094), .A1(n5757), .B0(n6111), .C0(n5996), .Y(n6109)
         );
  OAI21X4 U3669 ( .A0(n6079), .A1(n5664), .B0(n6080), .Y(n8182) );
  AOI211X4 U3670 ( .A0(n5095), .A1(n5667), .B0(n6081), .C0(n3364), .Y(n6079)
         );
  OAI21X4 U3671 ( .A0(n6133), .A1(n5826), .B0(n6134), .Y(n8200) );
  AOI211X4 U3672 ( .A0(n5094), .A1(n5829), .B0(n6135), .C0(n5996), .Y(n6133)
         );
  OAI21X4 U3673 ( .A0(n6103), .A1(n5736), .B0(n6104), .Y(n8190) );
  AOI211X4 U3674 ( .A0(n5094), .A1(n5739), .B0(n6105), .C0(n3364), .Y(n6103)
         );
  OAI21X4 U3675 ( .A0(n6145), .A1(n5862), .B0(n6146), .Y(n8204) );
  AOI211X4 U3676 ( .A0(n5094), .A1(n5865), .B0(n6147), .C0(n5996), .Y(n6145)
         );
  OAI21X4 U3677 ( .A0(n6112), .A1(n5763), .B0(n6113), .Y(n8193) );
  AOI211X4 U3678 ( .A0(n5094), .A1(n5766), .B0(n6114), .C0(n3364), .Y(n6112)
         );
  OAI21X4 U3679 ( .A0(n6097), .A1(n5718), .B0(n6098), .Y(n8188) );
  AOI211X4 U3680 ( .A0(n5095), .A1(n5721), .B0(n6099), .C0(n5996), .Y(n6097)
         );
  OAI21X4 U3681 ( .A0(n6124), .A1(n5799), .B0(n6125), .Y(n8197) );
  AOI211X4 U3682 ( .A0(n5094), .A1(n5802), .B0(n6126), .C0(n3364), .Y(n6124)
         );
  OAI21X4 U3683 ( .A0(n6106), .A1(n5745), .B0(n6107), .Y(n8191) );
  AOI211X4 U3684 ( .A0(n5094), .A1(n5748), .B0(n6108), .C0(n5996), .Y(n6106)
         );
  OAI21X4 U3685 ( .A0(n6139), .A1(n5844), .B0(n6140), .Y(n8202) );
  AOI211X4 U3686 ( .A0(n5094), .A1(n5847), .B0(n6141), .C0(n3364), .Y(n6139)
         );
  OAI21X4 U3687 ( .A0(n6043), .A1(n5556), .B0(n6044), .Y(n8170) );
  AOI211X4 U3688 ( .A0(n5095), .A1(n5559), .B0(n6045), .C0(n5996), .Y(n6043)
         );
  OAI21X4 U3689 ( .A0(n6121), .A1(n5790), .B0(n6122), .Y(n8196) );
  AOI211X4 U3690 ( .A0(n5094), .A1(n5793), .B0(n6123), .C0(n3364), .Y(n6121)
         );
  OAI21X4 U3691 ( .A0(n6118), .A1(n5781), .B0(n6119), .Y(n8195) );
  AOI211X4 U3692 ( .A0(n5094), .A1(n5784), .B0(n6120), .C0(n5996), .Y(n6118)
         );
  OAI21X4 U3693 ( .A0(n6142), .A1(n5853), .B0(n6143), .Y(n8203) );
  AOI211X4 U3694 ( .A0(n5094), .A1(n5856), .B0(n6144), .C0(n3364), .Y(n6142)
         );
  OAI21X4 U3695 ( .A0(n6130), .A1(n5817), .B0(n6131), .Y(n8199) );
  AOI211X4 U3696 ( .A0(n5094), .A1(n5820), .B0(n6132), .C0(n5996), .Y(n6130)
         );
  OAI21X4 U3697 ( .A0(n6115), .A1(n5772), .B0(n6116), .Y(n8194) );
  AOI211X4 U3698 ( .A0(n5094), .A1(n5775), .B0(n6117), .C0(n3364), .Y(n6115)
         );
  OAI21X4 U3699 ( .A0(n6148), .A1(n5871), .B0(n6149), .Y(n8205) );
  AOI211X4 U3700 ( .A0(n5094), .A1(n5874), .B0(n6150), .C0(n5996), .Y(n6148)
         );
  OAI21X4 U3701 ( .A0(n6007), .A1(n5448), .B0(n6008), .Y(n8158) );
  AOI211X4 U3702 ( .A0(n5096), .A1(n5451), .B0(n6009), .C0(n3364), .Y(n6007)
         );
  OAI21X4 U3703 ( .A0(n6013), .A1(n5466), .B0(n6014), .Y(n8160) );
  AOI211X4 U3704 ( .A0(n5096), .A1(n5469), .B0(n6015), .C0(n5996), .Y(n6013)
         );
  OAI21X4 U3705 ( .A0(n6082), .A1(n5673), .B0(n6083), .Y(n8183) );
  AOI211X4 U3706 ( .A0(n5095), .A1(n5676), .B0(n6084), .C0(n3364), .Y(n6082)
         );
  OAI21X4 U3707 ( .A0(n5998), .A1(n5421), .B0(n5999), .Y(n8155) );
  AOI211X4 U3708 ( .A0(n5096), .A1(n5424), .B0(n6000), .C0(n5996), .Y(n5998)
         );
  OAI21X4 U3709 ( .A0(n6004), .A1(n5439), .B0(n6005), .Y(n8157) );
  AOI211X4 U3710 ( .A0(n5096), .A1(n5442), .B0(n6006), .C0(n3364), .Y(n6004)
         );
  OAI21X4 U3711 ( .A0(n6067), .A1(n5628), .B0(n6068), .Y(n8178) );
  AOI211X4 U3712 ( .A0(n5095), .A1(n5631), .B0(n6069), .C0(n5996), .Y(n6067)
         );
  OAI21X4 U3713 ( .A0(n6073), .A1(n5646), .B0(n6074), .Y(n8180) );
  AOI211X4 U3714 ( .A0(n5095), .A1(n5649), .B0(n6075), .C0(n5996), .Y(n6073)
         );
  OAI21X4 U3715 ( .A0(n5992), .A1(n5408), .B0(n5993), .Y(n8154) );
  AOI211X4 U3716 ( .A0(n5096), .A1(n5412), .B0(n5995), .C0(n3364), .Y(n5992)
         );
  CLKBUFX20 U3717 ( .A(N2514), .Y(n3496) );
  OAI221X4 U3718 ( .A0(n5127), .A1(n3348), .B0(n5109), .B1(n8063), .C0(n8068), 
        .Y(N2514) );
  CLKINVX16 U3719 ( .A(n3481), .Y(n3482) );
  CLKINVX20 U3720 ( .A(n3481), .Y(n3484) );
  CLKINVX12 U3721 ( .A(n3481), .Y(n3485) );
  CLKINVX16 U3722 ( .A(n3481), .Y(n3483) );
  INVX16 U3723 ( .A(n3363), .Y(n3481) );
  AOI2BB2X2 U3724 ( .B0(n8065), .B1(n3751), .A0N(n3501), .A1N(n3523), .Y(n8070) );
  OR3X4 U3725 ( .A(n5350), .B(n5321), .C(n5379), .Y(n8087) );
  BUFX4 U3726 ( .A(n4123), .Y(n4130) );
  NAND4X6 U3727 ( .A(N2675), .B(N2674), .C(N2673), .D(n8088), .Y(n8080) );
  OAI222XL U3728 ( .A0(n5732), .A1(n5015), .B0(n5733), .B1(n5019), .C0(n5734), 
        .C1(n5023), .Y(n6892) );
  BUFX12 U3729 ( .A(N2486), .Y(n4947) );
  INVX4 U3730 ( .A(N2485), .Y(n5126) );
  OAI211X1 U3731 ( .A0(n5222), .A1(n5247), .B0(n5221), .C0(n5230), .Y(n5223)
         );
  INVX16 U3732 ( .A(n3488), .Y(n3489) );
  BUFX20 U3733 ( .A(n3737), .Y(n3742) );
  BUFX16 U3734 ( .A(n3921), .Y(n3931) );
  BUFX16 U3735 ( .A(n3520), .Y(n3522) );
  MX4XL U3736 ( .A(n4332), .B(n4330), .C(n4331), .D(n4329), .S0(n3503), .S1(
        n3495), .Y(n4333) );
  MX4X1 U3737 ( .A(n4230), .B(n4228), .C(n4229), .D(n4227), .S0(n5108), .S1(
        n3487), .Y(n4231) );
  MX4XL U3738 ( .A(n4397), .B(n4395), .C(n4396), .D(n4394), .S0(n3503), .S1(
        n3495), .Y(n4398) );
  BUFX16 U3739 ( .A(n3520), .Y(n3521) );
  BUFX20 U3740 ( .A(n3736), .Y(n3743) );
  MXI4X2 U3741 ( .A(n3957), .B(n3955), .C(n3956), .D(n3954), .S0(n4110), .S1(
        n3758), .Y(n3555) );
  MX4X1 U3742 ( .A(n4006), .B(n4004), .C(n4005), .D(n4003), .S0(n4108), .S1(
        n4135), .Y(n4007) );
  OAI32X1 U3743 ( .A0(n7945), .A1(n5053), .A2(n7940), .B0(n5065), .B1(n7931), 
        .Y(n7946) );
  OAI33X1 U3744 ( .A0(n7887), .A1(n5053), .A2(n7883), .B0(n7829), .B1(n7888), 
        .B2(n3562), .Y(n7889) );
  OAI33X1 U3745 ( .A0(n7788), .A1(n7196), .A2(n7784), .B0(n7730), .B1(n7789), 
        .B2(n3562), .Y(n7790) );
  OAI32X1 U3746 ( .A0(n7743), .A1(n7192), .A2(n7739), .B0(n5065), .B1(n3368), 
        .Y(n7742) );
  OAI32X1 U3747 ( .A0(n7743), .A1(n5053), .A2(n7739), .B0(n5065), .B1(n7730), 
        .Y(n7744) );
  OAI33X1 U3748 ( .A0(n7687), .A1(n7192), .A2(n7683), .B0(n4825), .B1(n7688), 
        .B2(n3562), .Y(n7686) );
  OAI33X1 U3749 ( .A0(n7687), .A1(n5053), .A2(n7683), .B0(n7629), .B1(n7688), 
        .B2(n5069), .Y(n7689) );
  OAI32X1 U3750 ( .A0(n7268), .A1(n5054), .A2(n7269), .B0(n3352), .B1(n7275), 
        .Y(n7276) );
  OAI33X1 U3751 ( .A0(n7272), .A1(n5053), .A2(n7268), .B0(n5069), .B1(n7273), 
        .B2(n7197), .Y(n7274) );
  OAI32X1 U3752 ( .A0(n7215), .A1(n5053), .A2(n7211), .B0(n7197), .B1(n5065), 
        .Y(n7216) );
  OAI32X1 U3753 ( .A0(n7211), .A1(n5054), .A2(n7212), .B0(n3352), .B1(n7218), 
        .Y(n7217) );
  OAI33X1 U3754 ( .A0(n8023), .A1(n5053), .A2(n8016), .B0(n7931), .B1(n8024), 
        .B2(n3558), .Y(n8026) );
  OAI32X1 U3755 ( .A0(n7971), .A1(n5053), .A2(n7965), .B0(n5067), .B1(n7931), 
        .Y(n7972) );
  OAI32X1 U3756 ( .A0(n7296), .A1(n5054), .A2(n7297), .B0(n3352), .B1(n7305), 
        .Y(n7306) );
  OAI33X1 U3757 ( .A0(n7300), .A1(n5053), .A2(n7296), .B0(n5071), .B1(n7301), 
        .B2(n7197), .Y(n7303) );
  OAI32X1 U3758 ( .A0(n7245), .A1(n5053), .A2(n7241), .B0(n7197), .B1(n5067), 
        .Y(n7246) );
  OAI32X1 U3759 ( .A0(n7241), .A1(n5054), .A2(n7242), .B0(n3351), .B1(n7248), 
        .Y(n7247) );
  OAI32X1 U3760 ( .A0(n7983), .A1(n5053), .A2(n7978), .B0(n5068), .B1(n7931), 
        .Y(n7984) );
  OAI33X1 U3761 ( .A0(n7927), .A1(n5053), .A2(n7920), .B0(n7931), .B1(n7929), 
        .B2(n5052), .Y(n7930) );
  OAI33X1 U3762 ( .A0(n7826), .A1(n5053), .A2(n7822), .B0(n7829), .B1(n7827), 
        .B2(n3548), .Y(n7828) );
  OAI33X1 U3763 ( .A0(n7727), .A1(n7192), .A2(n7723), .B0(n3368), .B1(n7728), 
        .B2(n5052), .Y(n7726) );
  OAI33X1 U3764 ( .A0(n7727), .A1(n5053), .A2(n7723), .B0(n7730), .B1(n7728), 
        .B2(n5052), .Y(n7729) );
  OAI33X1 U3765 ( .A0(n7625), .A1(n7192), .A2(n7621), .B0(n4825), .B1(n7627), 
        .B2(n5052), .Y(n7624) );
  OAI33X1 U3766 ( .A0(n7625), .A1(n5053), .A2(n7621), .B0(n7629), .B1(n7627), 
        .B2(n5052), .Y(n7628) );
  OAI33X1 U3767 ( .A0(n7525), .A1(n7192), .A2(n7521), .B0(n7526), .B1(n7527), 
        .B2(n5052), .Y(n7524) );
  OAI33X1 U3768 ( .A0(n7423), .A1(n5053), .A2(n7419), .B0(n7426), .B1(n7424), 
        .B2(n5052), .Y(n7425) );
  OAI32X1 U3769 ( .A0(n7318), .A1(n5054), .A2(n7319), .B0(n3351), .B1(n7327), 
        .Y(n7328) );
  OAI33X1 U3770 ( .A0(n7322), .A1(n5053), .A2(n7318), .B0(n7326), .B1(n7324), 
        .B2(n5052), .Y(n7325) );
  OAI32X1 U3771 ( .A0(n7260), .A1(n5051), .A2(n7256), .B0(n7193), .B1(n5068), 
        .Y(n7259) );
  OAI32X1 U3772 ( .A0(n7260), .A1(n5053), .A2(n7256), .B0(n7197), .B1(n5068), 
        .Y(n7261) );
  OAI32X1 U3773 ( .A0(n7256), .A1(n5054), .A2(n7257), .B0(n3352), .B1(n7263), 
        .Y(n7262) );
  OAI33X1 U3774 ( .A0(n7957), .A1(n7192), .A2(n7952), .B0(n7928), .B1(n7958), 
        .B2(n5066), .Y(n7956) );
  OAI33X1 U3775 ( .A0(n7957), .A1(n5053), .A2(n7952), .B0(n7931), .B1(n7958), 
        .B2(n5066), .Y(n7959) );
  OAI32X1 U3776 ( .A0(n7952), .A1(n5059), .A2(n7953), .B0(n3351), .B1(n7960), 
        .Y(n7961) );
  OAI33X1 U3777 ( .A0(n7853), .A1(n5053), .A2(n7849), .B0(n7829), .B1(n7854), 
        .B2(n5066), .Y(n7855) );
  OAI32X1 U3778 ( .A0(n7800), .A1(n5053), .A2(n7796), .B0(n5070), .B1(n7730), 
        .Y(n7801) );
  OAI33X1 U3779 ( .A0(n7754), .A1(n7192), .A2(n7750), .B0(n3368), .B1(n7755), 
        .B2(n3561), .Y(n7753) );
  OAI33X1 U3780 ( .A0(n7754), .A1(n5053), .A2(n7750), .B0(n7730), .B1(n7755), 
        .B2(n5066), .Y(n7756) );
  OAI33X1 U3781 ( .A0(n7653), .A1(n7192), .A2(n7649), .B0(n4825), .B1(n7654), 
        .B2(n5066), .Y(n7652) );
  OAI33X1 U3782 ( .A0(n7653), .A1(n5053), .A2(n7649), .B0(n7629), .B1(n7654), 
        .B2(n3561), .Y(n7655) );
  OAI33X1 U3783 ( .A0(n7553), .A1(n7192), .A2(n7549), .B0(n7526), .B1(n7554), 
        .B2(n5066), .Y(n7552) );
  OAI33X1 U3784 ( .A0(n7450), .A1(n5053), .A2(n7446), .B0(n7426), .B1(n7451), 
        .B2(n5066), .Y(n7452) );
  OAI32X1 U3785 ( .A0(n7346), .A1(n5054), .A2(n7347), .B0(n3351), .B1(n7353), 
        .Y(n7354) );
  OAI33X1 U3786 ( .A0(n7350), .A1(n5053), .A2(n7346), .B0(n7326), .B1(n7351), 
        .B2(n3561), .Y(n7352) );
  OAI32X1 U3787 ( .A0(n7287), .A1(n7192), .A2(n7283), .B0(n7193), .B1(n5070), 
        .Y(n7286) );
  OAI32X1 U3788 ( .A0(n7287), .A1(n5053), .A2(n7283), .B0(n7197), .B1(n5070), 
        .Y(n7288) );
  OAI32X1 U3789 ( .A0(n7283), .A1(n5054), .A2(n7284), .B0(n3351), .B1(n7290), 
        .Y(n7289) );
  AOI2BB2XL U3790 ( .B0(n8079), .B1(n4947), .A0N(n7308), .A1N(n8080), .Y(n8078) );
  AOI2BB2XL U3791 ( .B0(n8079), .B1(n5125), .A0N(n7307), .A1N(n8080), .Y(n8081) );
  MX4XL U3792 ( .A(n4041), .B(n4039), .C(n4040), .D(n4038), .S0(n4108), .S1(
        n4135), .Y(n4042) );
  AOI2BB2XL U3793 ( .B0(n8065), .B1(n4947), .A0N(n7308), .A1N(n3523), .Y(n8064) );
  OAI33X1 U3794 ( .A0(n7229), .A1(n7192), .A2(n7225), .B0(n5066), .B1(n7230), 
        .B2(n7193), .Y(n7228) );
  OAI32X1 U3795 ( .A0(n7225), .A1(n5054), .A2(n7226), .B0(n3351), .B1(n7232), 
        .Y(n7233) );
  OAI33X1 U3796 ( .A0(n7229), .A1(n5053), .A2(n7225), .B0(n5066), .B1(n7230), 
        .B2(n7197), .Y(n7231) );
  OAI222XL U3797 ( .A0(n5768), .A1(n5015), .B0(n5769), .B1(n5018), .C0(n5770), 
        .C1(n5023), .Y(n6904) );
  INVX3 U3798 ( .A(n7993), .Y(n5968) );
  CLKINVX1 U3799 ( .A(n7947), .Y(n5930) );
  CLKINVX1 U3800 ( .A(n7886), .Y(n5896) );
  CLKINVX1 U3801 ( .A(n7889), .Y(n5895) );
  CLKINVX1 U3802 ( .A(n7787), .Y(n5824) );
  CLKINVX1 U3803 ( .A(n7790), .Y(n5823) );
  CLKINVX1 U3804 ( .A(n7742), .Y(n5788) );
  CLKINVX1 U3805 ( .A(n7686), .Y(n5752) );
  CLKINVX1 U3806 ( .A(n7689), .Y(n5751) );
  NAND2X2 U3807 ( .A(n5042), .B(n4914), .Y(n5745) );
  INVX3 U3808 ( .A(n7641), .Y(n5716) );
  OAI32X1 U3809 ( .A0(n7642), .A1(n7196), .A2(n7638), .B0(n5065), .B1(n7629), 
        .Y(n7643) );
  INVX3 U3810 ( .A(n7591), .Y(n5678) );
  CLKINVX1 U3811 ( .A(n7589), .Y(n5679) );
  NAND2X2 U3812 ( .A(n5041), .B(n4901), .Y(n5637) );
  CLKINVX1 U3813 ( .A(n7271), .Y(n5464) );
  INVX1 U3814 ( .A(n8022), .Y(n5991) );
  CLKINVX1 U3815 ( .A(n8032), .Y(n5989) );
  OAI22XL U3816 ( .A0(n7293), .A1(n7918), .B0(n8012), .B1(n3344), .Y(n5981) );
  OAI22XL U3817 ( .A0(n7238), .A1(n7918), .B0(n7964), .B1(n3344), .Y(n5945) );
  OAI33X1 U3818 ( .A0(n7910), .A1(n7192), .A2(n7906), .B0(n3369), .B1(n7911), 
        .B2(n3558), .Y(n7909) );
  OAI22XL U3819 ( .A0(n7293), .A1(n7819), .B0(n7905), .B1(n3344), .Y(n5909) );
  OAI22XL U3820 ( .A0(n7238), .A1(n7819), .B0(n7860), .B1(n3344), .Y(n5873) );
  OAI33X1 U3821 ( .A0(n7811), .A1(n5053), .A2(n7807), .B0(n7730), .B1(n7812), 
        .B2(n5071), .Y(n7814) );
  INVX3 U3822 ( .A(n7664), .Y(n5734) );
  OAI32X1 U3823 ( .A0(n7665), .A1(n7196), .A2(n7661), .B0(n3549), .B1(n7629), 
        .Y(n7666) );
  OAI22XL U3824 ( .A0(n7293), .A1(n7518), .B0(n7605), .B1(n3344), .Y(n5693) );
  OAI22XL U3825 ( .A0(n7238), .A1(n7518), .B0(n7560), .B1(n3344), .Y(n5657) );
  OAI22XL U3826 ( .A0(n7293), .A1(n7416), .B0(n7502), .B1(n3344), .Y(n5621) );
  OAI22XL U3827 ( .A0(n7238), .A1(n7416), .B0(n7457), .B1(n3344), .Y(n5585) );
  OAI33X1 U3828 ( .A0(n7408), .A1(n5053), .A2(n7403), .B0(n7326), .B1(n7409), 
        .B2(n5071), .Y(n7411) );
  OAI22XL U3829 ( .A0(n7293), .A1(n7314), .B0(n7402), .B1(n3344), .Y(n5549) );
  INVX3 U3830 ( .A(n7364), .Y(n5516) );
  OAI32X1 U3831 ( .A0(n7358), .A1(n5054), .A2(n7359), .B0(n3352), .B1(n7365), 
        .Y(n7364) );
  CLKINVX1 U3832 ( .A(n7299), .Y(n5482) );
  OAI22XL U3833 ( .A0(n7253), .A1(n7918), .B0(n7977), .B1(n3344), .Y(n5954) );
  CLKINVX1 U3834 ( .A(n7926), .Y(n5923) );
  OAI32X1 U3835 ( .A0(n7872), .A1(n5058), .A2(n7873), .B0(n3352), .B1(n7879), 
        .Y(n7878) );
  OAI22XL U3836 ( .A0(n7253), .A1(n7819), .B0(n7871), .B1(n3344), .Y(n5882) );
  CLKINVX1 U3837 ( .A(n7825), .Y(n5851) );
  CLKINVX1 U3838 ( .A(n7828), .Y(n5850) );
  OAI32XL U3839 ( .A0(n7777), .A1(n7192), .A2(n7773), .B0(n5068), .B1(n3368), 
        .Y(n7776) );
  OAI22XL U3840 ( .A0(n7253), .A1(n7720), .B0(n7772), .B1(n3344), .Y(n5810) );
  CLKINVX1 U3841 ( .A(n7726), .Y(n5779) );
  CLKINVX1 U3842 ( .A(n7729), .Y(n5778) );
  CLKINVX1 U3843 ( .A(n7624), .Y(n5707) );
  CLKINVX1 U3844 ( .A(n7528), .Y(n5634) );
  OAI22XL U3845 ( .A0(n7253), .A1(n7416), .B0(n7468), .B1(n3344), .Y(n5594) );
  INVX3 U3846 ( .A(n7428), .Y(n5561) );
  CLKINVX1 U3847 ( .A(n7422), .Y(n5563) );
  INVX3 U3848 ( .A(n7375), .Y(n5525) );
  OAI32X1 U3849 ( .A0(n7369), .A1(n5054), .A2(n7370), .B0(n3352), .B1(n7376), 
        .Y(n7375) );
  CLKINVX1 U3850 ( .A(n7321), .Y(n5491) );
  INVX3 U3851 ( .A(n7199), .Y(n5415) );
  CLKINVX1 U3852 ( .A(n7961), .Y(n5939) );
  OAI32X1 U3853 ( .A0(n7895), .A1(n5058), .A2(n7896), .B0(n3352), .B1(n7902), 
        .Y(n7901) );
  CLKINVX1 U3854 ( .A(n7852), .Y(n5869) );
  CLKINVX1 U3855 ( .A(n7799), .Y(n5833) );
  CLKINVX1 U3856 ( .A(n7753), .Y(n5797) );
  CLKINVX1 U3857 ( .A(n7756), .Y(n5796) );
  INVX3 U3858 ( .A(n7698), .Y(n5761) );
  NAND2X2 U3859 ( .A(n5042), .B(n4915), .Y(n5754) );
  CLKINVX1 U3860 ( .A(n7652), .Y(n5725) );
  CLKINVX1 U3861 ( .A(n7555), .Y(n5652) );
  NAND2X2 U3862 ( .A(n5042), .B(n4902), .Y(n5646) );
  INVX3 U3863 ( .A(n7454), .Y(n5579) );
  CLKINVX1 U3864 ( .A(n7449), .Y(n5581) );
  CLKINVX1 U3865 ( .A(n7349), .Y(n5509) );
  CLKINVX1 U3866 ( .A(n7352), .Y(n5508) );
  INVX12 U3867 ( .A(n5078), .Y(n5077) );
  CLKINVX1 U3868 ( .A(n7228), .Y(n5437) );
  CLKINVX1 U3869 ( .A(n7231), .Y(n5436) );
  NOR2BX1 U3870 ( .AN(N2773), .B(N2781), .Y(n5191) );
  NAND2BX1 U3871 ( .AN(n3944), .B(N2779), .Y(n5171) );
  NOR2X1 U3872 ( .A(n5162), .B(n5174), .Y(n5175) );
  NAND2BX1 U3873 ( .AN(n5184), .B(n5166), .Y(n5179) );
  AND2X2 U3874 ( .A(n5193), .B(n5203), .Y(n5200) );
  NOR2X1 U3875 ( .A(n5194), .B(n5206), .Y(n5207) );
  CLKINVX1 U3876 ( .A(n5135), .Y(n5158) );
  NOR2X1 U3877 ( .A(n5157), .B(n4867), .Y(n5154) );
  AOI211X1 U3878 ( .A0(n5285), .A1(n5297), .B0(n5284), .C0(n5300), .Y(n5286)
         );
  AOI31X1 U3879 ( .A0(n5298), .A1(n5283), .A2(n5282), .B0(n5295), .Y(n5285) );
  AOI211X1 U3880 ( .A0(n5375), .A1(n5387), .B0(n5374), .C0(n5390), .Y(n5376)
         );
  AOI31X1 U3881 ( .A0(n5331), .A1(n5330), .A2(n5329), .B0(n5328), .Y(n5335) );
  NAND3BX1 U3882 ( .AN(n5327), .B(n5326), .C(n5325), .Y(n5331) );
  OAI211X1 U3883 ( .A0(n5077), .A1(n5324), .B0(n5323), .C0(n5322), .Y(n5326)
         );
  AOI31X1 U3884 ( .A0(n5360), .A1(n5359), .A2(n5358), .B0(n5357), .Y(n5364) );
  NAND3BX1 U3885 ( .AN(n5356), .B(n5355), .C(n5354), .Y(n5360) );
  OAI211X1 U3886 ( .A0(n5077), .A1(n5353), .B0(n5352), .C0(n5351), .Y(n5355)
         );
  CLKINVX1 U3887 ( .A(n3541), .Y(n5264) );
  OA21XL U3888 ( .A0(n4873), .A1(n5261), .B0(n5260), .Y(n3433) );
  CLKBUFX3 U3889 ( .A(n5345), .Y(n3492) );
  NAND2BX1 U3890 ( .AN(n5245), .B(n5228), .Y(n5240) );
  NOR2X1 U3891 ( .A(n5250), .B(n4861), .Y(n5246) );
  NOR2X1 U3892 ( .A(n5188), .B(n5101), .Y(n5185) );
  NAND2X1 U3893 ( .A(n4867), .B(n5157), .Y(n5151) );
  NOR2X2 U3894 ( .A(n5219), .B(N2767), .Y(n5216) );
  MX4X1 U3895 ( .A(n4145), .B(n4143), .C(n4144), .D(n4142), .S0(n5108), .S1(
        n3487), .Y(n4146) );
  MX4X1 U3896 ( .A(\ImageBuffer[20][2] ), .B(\ImageBuffer[21][2] ), .C(
        \ImageBuffer[22][2] ), .D(\ImageBuffer[23][2] ), .S0(n3513), .S1(n3471), .Y(n4371) );
  CLKINVX4 U3897 ( .A(n3940), .Y(n3488) );
  NAND2X2 U3898 ( .A(cmd[3]), .B(n3476), .Y(n8029) );
  BUFX4 U3899 ( .A(n5113), .Y(n4316) );
  MX4X1 U3900 ( .A(\ImageBuffer[60][1] ), .B(\ImageBuffer[61][1] ), .C(
        \ImageBuffer[62][1] ), .D(\ImageBuffer[63][1] ), .S0(n3939), .S1(n4311), .Y(n4157) );
  MX4X1 U3901 ( .A(\ImageBuffer[48][1] ), .B(\ImageBuffer[49][1] ), .C(
        \ImageBuffer[50][1] ), .D(\ImageBuffer[51][1] ), .S0(n3939), .S1(n4317), .Y(n4160) );
  MX4X1 U3902 ( .A(\ImageBuffer[56][1] ), .B(\ImageBuffer[57][1] ), .C(
        \ImageBuffer[58][1] ), .D(\ImageBuffer[59][1] ), .S0(n3497), .S1(n4306), .Y(n4158) );
  MX4X1 U3903 ( .A(\ImageBuffer[36][1] ), .B(\ImageBuffer[37][1] ), .C(
        \ImageBuffer[38][1] ), .D(\ImageBuffer[39][1] ), .S0(n3939), .S1(n4314), .Y(n4164) );
  MX4X1 U3904 ( .A(\ImageBuffer[44][1] ), .B(\ImageBuffer[45][1] ), .C(
        \ImageBuffer[46][1] ), .D(\ImageBuffer[47][1] ), .S0(n3939), .S1(n4305), .Y(n4162) );
  MX4X1 U3905 ( .A(n3981), .B(n3979), .C(n3980), .D(n3978), .S0(n4108), .S1(
        n4135), .Y(n3982) );
  CLKBUFX3 U3906 ( .A(n3945), .Y(N2786) );
  CLKBUFX3 U3907 ( .A(N2505), .Y(n3520) );
  CLKBUFX3 U3908 ( .A(n3745), .Y(n3736) );
  NAND3BX1 U3909 ( .AN(n5295), .B(n5294), .C(n5293), .Y(n5299) );
  MX4X1 U3910 ( .A(n3773), .B(n3771), .C(n3772), .D(n3770), .S0(n3934), .S1(
        n3409), .Y(n3774) );
  MX4X1 U3911 ( .A(n3966), .B(n3964), .C(n3965), .D(n3963), .S0(n4109), .S1(
        n3758), .Y(n3967) );
  MX4X1 U3912 ( .A(\ImageBuffer[8][0] ), .B(\ImageBuffer[9][0] ), .C(
        \ImageBuffer[10][0] ), .D(\ImageBuffer[11][0] ), .S0(n3735), .S1(n4132), .Y(n3964) );
  MX4X1 U3913 ( .A(\ImageBuffer[0][0] ), .B(\ImageBuffer[1][0] ), .C(
        \ImageBuffer[2][0] ), .D(\ImageBuffer[3][0] ), .S0(n3735), .S1(n4126), 
        .Y(n3966) );
  CLKINVX1 U3914 ( .A(n3962), .Y(n3554) );
  MX4X1 U3915 ( .A(n3961), .B(n3959), .C(n3960), .D(n3958), .S0(n4108), .S1(
        n3758), .Y(n3962) );
  MX4X1 U3916 ( .A(\ImageBuffer[28][0] ), .B(\ImageBuffer[29][0] ), .C(
        \ImageBuffer[30][0] ), .D(\ImageBuffer[31][0] ), .S0(n4114), .S1(n3749), .Y(n3958) );
  MX4X1 U3917 ( .A(\ImageBuffer[20][0] ), .B(\ImageBuffer[21][0] ), .C(
        \ImageBuffer[22][0] ), .D(\ImageBuffer[23][0] ), .S0(n4114), .S1(n3749), .Y(n3960) );
  MX4X1 U3918 ( .A(\ImageBuffer[4][2] ), .B(\ImageBuffer[5][2] ), .C(
        \ImageBuffer[6][2] ), .D(\ImageBuffer[7][2] ), .S0(n3515), .S1(n3471), 
        .Y(n4376) );
  MX4X1 U3919 ( .A(\ImageBuffer[12][2] ), .B(\ImageBuffer[13][2] ), .C(
        \ImageBuffer[14][2] ), .D(\ImageBuffer[15][2] ), .S0(n3516), .S1(n3471), .Y(n4374) );
  MX4X1 U3920 ( .A(\ImageBuffer[8][2] ), .B(\ImageBuffer[9][2] ), .C(
        \ImageBuffer[10][2] ), .D(\ImageBuffer[11][2] ), .S0(n3511), .S1(n3472), .Y(n4375) );
  MX4X1 U3921 ( .A(\ImageBuffer[0][2] ), .B(\ImageBuffer[1][2] ), .C(
        \ImageBuffer[2][2] ), .D(\ImageBuffer[3][2] ), .S0(n3512), .S1(n3473), 
        .Y(n4377) );
  MX4X1 U3922 ( .A(\ImageBuffer[48][2] ), .B(\ImageBuffer[49][2] ), .C(
        \ImageBuffer[50][2] ), .D(\ImageBuffer[51][2] ), .S0(n3515), .S1(n3472), .Y(n4362) );
  MX4X1 U3923 ( .A(\ImageBuffer[56][2] ), .B(\ImageBuffer[57][2] ), .C(
        \ImageBuffer[58][2] ), .D(\ImageBuffer[59][2] ), .S0(n3517), .S1(n3473), .Y(n4360) );
  MX4X1 U3924 ( .A(\ImageBuffer[52][2] ), .B(\ImageBuffer[53][2] ), .C(
        \ImageBuffer[54][2] ), .D(\ImageBuffer[55][2] ), .S0(n3513), .S1(n3472), .Y(n4361) );
  MX4X1 U3925 ( .A(\ImageBuffer[60][2] ), .B(\ImageBuffer[61][2] ), .C(
        \ImageBuffer[62][2] ), .D(\ImageBuffer[63][2] ), .S0(n3514), .S1(n3473), .Y(n4359) );
  MX4X1 U3926 ( .A(\ImageBuffer[44][2] ), .B(\ImageBuffer[45][2] ), .C(
        \ImageBuffer[46][2] ), .D(\ImageBuffer[47][2] ), .S0(n3516), .S1(n3472), .Y(n4364) );
  MX4X1 U3927 ( .A(\ImageBuffer[32][2] ), .B(\ImageBuffer[33][2] ), .C(
        \ImageBuffer[34][2] ), .D(\ImageBuffer[35][2] ), .S0(n3513), .S1(n3474), .Y(n4367) );
  MX4X1 U3928 ( .A(\ImageBuffer[36][2] ), .B(\ImageBuffer[37][2] ), .C(
        \ImageBuffer[38][2] ), .D(\ImageBuffer[39][2] ), .S0(n3511), .S1(n3471), .Y(n4366) );
  MX4X1 U3929 ( .A(\ImageBuffer[40][2] ), .B(\ImageBuffer[41][2] ), .C(
        \ImageBuffer[42][2] ), .D(\ImageBuffer[43][2] ), .S0(n3512), .S1(n3474), .Y(n4365) );
  MX4X1 U3930 ( .A(n4372), .B(n4370), .C(n4371), .D(n4369), .S0(n3503), .S1(
        n3495), .Y(n4373) );
  MX4X1 U3931 ( .A(\ImageBuffer[28][2] ), .B(\ImageBuffer[29][2] ), .C(
        \ImageBuffer[30][2] ), .D(\ImageBuffer[31][2] ), .S0(n3514), .S1(n3472), .Y(n4369) );
  MX4X1 U3932 ( .A(\ImageBuffer[16][2] ), .B(\ImageBuffer[17][2] ), .C(
        \ImageBuffer[18][2] ), .D(\ImageBuffer[19][2] ), .S0(n3514), .S1(n3473), .Y(n4372) );
  MX4X1 U3933 ( .A(\ImageBuffer[24][2] ), .B(\ImageBuffer[25][2] ), .C(
        \ImageBuffer[26][2] ), .D(\ImageBuffer[27][2] ), .S0(n3513), .S1(n3474), .Y(n4370) );
  MX4X1 U3934 ( .A(n3991), .B(n3989), .C(n3990), .D(n3988), .S0(n4108), .S1(
        n4135), .Y(n3992) );
  MX4X1 U3935 ( .A(n3996), .B(n3994), .C(n3995), .D(n3993), .S0(n4108), .S1(
        n4135), .Y(n3997) );
  MX4X1 U3936 ( .A(\ImageBuffer[0][3] ), .B(\ImageBuffer[1][3] ), .C(
        \ImageBuffer[2][3] ), .D(\ImageBuffer[3][3] ), .S0(n3742), .S1(n4133), 
        .Y(n3651) );
  MX4X1 U3937 ( .A(n3636), .B(n3634), .C(n3635), .D(n3633), .S0(n3734), .S1(
        n3758), .Y(n3637) );
  MX4X1 U3938 ( .A(n3783), .B(n3781), .C(n3782), .D(n3780), .S0(n3934), .S1(
        n3409), .Y(n3784) );
  XOR2X1 U3939 ( .A(N2495), .B(n3470), .Y(N2501) );
  MX4X1 U3940 ( .A(n3858), .B(n3856), .C(n3857), .D(n3855), .S0(n3933), .S1(
        n3409), .Y(n3859) );
  MX4X1 U3941 ( .A(\ImageBuffer[4][5] ), .B(\ImageBuffer[5][5] ), .C(
        \ImageBuffer[6][5] ), .D(\ImageBuffer[7][5] ), .S0(n3743), .S1(n4123), 
        .Y(n3690) );
  MX4X1 U3942 ( .A(\ImageBuffer[20][5] ), .B(\ImageBuffer[21][5] ), .C(
        \ImageBuffer[22][5] ), .D(\ImageBuffer[23][5] ), .S0(n3743), .S1(n4131), .Y(n3685) );
  MX4X1 U3943 ( .A(\ImageBuffer[24][5] ), .B(\ImageBuffer[25][5] ), .C(
        \ImageBuffer[26][5] ), .D(\ImageBuffer[27][5] ), .S0(n3743), .S1(n3754), .Y(n3684) );
  MX4X1 U3944 ( .A(n4342), .B(n4340), .C(n4341), .D(n4339), .S0(n3503), .S1(
        n3495), .Y(n4343) );
  INVX16 U3945 ( .A(n3504), .Y(n3473) );
  INVX16 U3946 ( .A(n3504), .Y(n3471) );
  MX4X1 U3947 ( .A(n4046), .B(n4044), .C(n4045), .D(n4043), .S0(n4109), .S1(
        n4136), .Y(n4047) );
  CLKBUFX8 U3948 ( .A(n3748), .Y(n3753) );
  MX4X1 U3949 ( .A(n4612), .B(n4610), .C(n4611), .D(n4609), .S0(n3496), .S1(
        n4640), .Y(n4613) );
  MX4X1 U3950 ( .A(\ImageBuffer[36][6] ), .B(\ImageBuffer[37][6] ), .C(
        \ImageBuffer[38][6] ), .D(\ImageBuffer[39][6] ), .S0(n4118), .S1(n4128), .Y(n4075) );
  MX4X1 U3951 ( .A(\ImageBuffer[20][6] ), .B(\ImageBuffer[21][6] ), .C(
        \ImageBuffer[22][6] ), .D(\ImageBuffer[23][6] ), .S0(n4118), .S1(n3754), .Y(n4080) );
  MX4X1 U3952 ( .A(\ImageBuffer[28][6] ), .B(\ImageBuffer[29][6] ), .C(
        \ImageBuffer[30][6] ), .D(\ImageBuffer[31][6] ), .S0(n4118), .S1(n4133), .Y(n4078) );
  INVX16 U3953 ( .A(n3502), .Y(n3503) );
  INVX8 U3954 ( .A(n3494), .Y(n3495) );
  MX4X1 U3955 ( .A(n4492), .B(n4490), .C(n4491), .D(n4489), .S0(n3496), .S1(
        n4641), .Y(n4493) );
  MX4X1 U3956 ( .A(n4337), .B(n4335), .C(n4336), .D(n4334), .S0(n3503), .S1(
        n3495), .Y(n4338) );
  MX4X1 U3957 ( .A(n4327), .B(n4325), .C(n4326), .D(n4324), .S0(n3503), .S1(
        n3495), .Y(n4328) );
  MX4X1 U3958 ( .A(n4378), .B(n4368), .C(n4373), .D(n4363), .S0(N2510), .S1(
        N2509), .Y(N2747) );
  MX4X1 U3959 ( .A(n4367), .B(n4365), .C(n4366), .D(n4364), .S0(n3503), .S1(
        n3495), .Y(n4368) );
  MX4X1 U3960 ( .A(n4362), .B(n4360), .C(n4361), .D(n4359), .S0(n3503), .S1(
        n3495), .Y(n4363) );
  MX4X1 U3961 ( .A(n4377), .B(n4375), .C(n4376), .D(n4374), .S0(n3503), .S1(
        n3495), .Y(n4378) );
  MX4X1 U3962 ( .A(n4537), .B(n4535), .C(n4536), .D(n4534), .S0(n3496), .S1(
        n4639), .Y(n4538) );
  MX4X1 U3963 ( .A(n4522), .B(n4520), .C(n4521), .D(n4519), .S0(n3496), .S1(
        n4639), .Y(n4523) );
  CLKINVX1 U3964 ( .A(n7994), .Y(n7991) );
  CLKINVX1 U3965 ( .A(n7945), .Y(n7941) );
  CLKINVX1 U3966 ( .A(n7887), .Y(n7884) );
  CLKINVX1 U3967 ( .A(n7788), .Y(n7785) );
  CLKINVX1 U3968 ( .A(n7743), .Y(n7740) );
  CLKINVX1 U3969 ( .A(n7687), .Y(n7684) );
  CLKINVX1 U3970 ( .A(n7642), .Y(n7639) );
  OAI32X1 U3971 ( .A0(n7480), .A1(n5055), .A2(n7481), .B0(n3351), .B1(n7487), 
        .Y(n7488) );
  OAI33X1 U3972 ( .A0(n7484), .A1(n7192), .A2(n7480), .B0(n3367), .B1(n7485), 
        .B2(n5069), .Y(n7483) );
  OAI33X1 U3973 ( .A0(n7484), .A1(n5053), .A2(n7480), .B0(n7426), .B1(n7485), 
        .B2(n5069), .Y(n7486) );
  OAI32X1 U3974 ( .A0(n7380), .A1(n5055), .A2(n7381), .B0(n3351), .B1(n7387), 
        .Y(n7388) );
  OAI33X1 U3975 ( .A0(n7384), .A1(n5053), .A2(n7380), .B0(n7326), .B1(n7385), 
        .B2(n5069), .Y(n7386) );
  CLKINVX1 U3976 ( .A(n7910), .Y(n7907) );
  OAI32X1 U3977 ( .A0(n7766), .A1(n5053), .A2(n7762), .B0(n3549), .B1(n7730), 
        .Y(n7767) );
  CLKINVX1 U3978 ( .A(n7766), .Y(n7763) );
  CLKINVX1 U3979 ( .A(n7711), .Y(n7707) );
  CLKINVX1 U3980 ( .A(n7665), .Y(n7662) );
  CLKINVX1 U3981 ( .A(n7983), .Y(n7979) );
  CLKINVX1 U3982 ( .A(n7927), .Y(n7921) );
  CLKINVX1 U3983 ( .A(n7876), .Y(n7873) );
  CLKINVX1 U3984 ( .A(n7826), .Y(n7823) );
  CLKINVX1 U3985 ( .A(n7777), .Y(n7774) );
  CLKINVX1 U3986 ( .A(n7727), .Y(n7724) );
  CLKINVX1 U3987 ( .A(n7676), .Y(n7673) );
  CLKINVX1 U3988 ( .A(n7625), .Y(n7622) );
  CLKINVX1 U3989 ( .A(n8006), .Y(n8003) );
  CLKINVX1 U3990 ( .A(n7957), .Y(n7953) );
  CLKINVX1 U3991 ( .A(n7899), .Y(n7896) );
  CLKINVX1 U3992 ( .A(n7853), .Y(n7850) );
  CLKINVX1 U3993 ( .A(n7800), .Y(n7797) );
  BUFX4 U3994 ( .A(N2760), .Y(n4869) );
  CLKINVX1 U3995 ( .A(n7754), .Y(n7751) );
  MX4X1 U3996 ( .A(n3611), .B(n3609), .C(n3610), .D(n3608), .S0(n3734), .S1(
        n3758), .Y(n3612) );
  BUFX6 U3997 ( .A(N2764), .Y(n4873) );
  MX4X2 U3998 ( .A(n3799), .B(n3789), .C(n3794), .D(n3784), .S0(N2492), .S1(
        N2491), .Y(N2764) );
  MX4X1 U3999 ( .A(n3798), .B(n3796), .C(n3797), .D(n3795), .S0(n3933), .S1(
        n3409), .Y(n3799) );
  MX4X2 U4000 ( .A(n3788), .B(n3786), .C(n3787), .D(n3785), .S0(n3934), .S1(
        n3409), .Y(n3789) );
  MX4X1 U4001 ( .A(n3656), .B(n3654), .C(n3655), .D(n3653), .S0(n3734), .S1(
        n3758), .Y(n3657) );
  CLKBUFX3 U4002 ( .A(n7626), .Y(n4825) );
  CLKINVX1 U4003 ( .A(n7699), .Y(n7696) );
  CLKINVX1 U4004 ( .A(n7653), .Y(n7650) );
  MX4X1 U4005 ( .A(n4235), .B(n4233), .C(n4234), .D(n4232), .S0(n5108), .S1(
        n3487), .Y(n4236) );
  MX4X1 U4006 ( .A(n4220), .B(n4218), .C(n4219), .D(n4217), .S0(n5108), .S1(
        n3487), .Y(n4221) );
  MX4X1 U4007 ( .A(n4225), .B(n4223), .C(n4224), .D(n4222), .S0(n5108), .S1(
        n3487), .Y(n4226) );
  MX4X2 U4008 ( .A(n4216), .B(n4206), .C(n4211), .D(n4201), .S0(N2504), .S1(
        N2503), .Y(N2770) );
  MX4X1 U4009 ( .A(n4387), .B(n4385), .C(n4386), .D(n4384), .S0(n3503), .S1(
        n3495), .Y(n4388) );
  MX4X1 U4010 ( .A(n4392), .B(n4390), .C(n4391), .D(n4389), .S0(n3503), .S1(
        n3495), .Y(n4393) );
  MX4X1 U4011 ( .A(n4572), .B(n4570), .C(n4571), .D(n4569), .S0(n3496), .S1(
        n4639), .Y(n4573) );
  MX4X1 U4012 ( .A(n4562), .B(n4560), .C(n4561), .D(n4559), .S0(n3496), .S1(
        n4639), .Y(n4563) );
  MX4X1 U4013 ( .A(n4407), .B(n4405), .C(n4406), .D(n4404), .S0(n3503), .S1(
        n3495), .Y(n4408) );
  MX4X1 U4014 ( .A(n4402), .B(n4400), .C(n4401), .D(n4399), .S0(n3503), .S1(
        n3495), .Y(n4403) );
  MX4X1 U4015 ( .A(n4438), .B(n4428), .C(n4433), .D(n4423), .S0(N2510), .S1(
        N2509), .Y(N2744) );
  MX4X1 U4016 ( .A(n4437), .B(n4435), .C(n4436), .D(n4434), .S0(n3503), .S1(
        n3495), .Y(n4438) );
  NAND2X1 U4017 ( .A(sum[8]), .B(n5987), .Y(n3567) );
  MX4X1 U4018 ( .A(n4632), .B(n4630), .C(n4631), .D(n4629), .S0(n3496), .S1(
        n4640), .Y(n4633) );
  INVX3 U4019 ( .A(N2493), .Y(n5121) );
  CLKINVX1 U4020 ( .A(n8620), .Y(n7968) );
  INVX16 U4021 ( .A(N2494), .Y(n5117) );
  BUFX8 U4022 ( .A(n4134), .Y(n4123) );
  CLKXOR2X4 U4023 ( .A(\r2549/carry[5] ), .B(n4947), .Y(N2492) );
  NAND2X1 U4024 ( .A(N2757), .B(n5988), .Y(n3442) );
  NAND2X1 U4025 ( .A(sum[4]), .B(n5987), .Y(n3543) );
  NAND2X1 U4026 ( .A(N2747), .B(n4943), .Y(n3542) );
  CLKINVX1 U4027 ( .A(n7765), .Y(n5806) );
  OAI22XL U4028 ( .A0(n7238), .A1(n7720), .B0(n7761), .B1(n3344), .Y(n5801) );
  INVX12 U4029 ( .A(n6187), .Y(n3364) );
  INVX12 U4030 ( .A(n6583), .Y(n6390) );
  MX4X1 U4031 ( .A(n4418), .B(n4408), .C(n4413), .D(n4403), .S0(N2510), .S1(
        N2509), .Y(N2745) );
  CLKBUFX8 U4032 ( .A(n3947), .Y(n5093) );
  INVX12 U4033 ( .A(n3469), .Y(n6192) );
  MX4X1 U4034 ( .A(n4598), .B(n4588), .C(n4593), .D(n4583), .S0(N2516), .S1(
        N2515), .Y(N2752) );
  INVX12 U4035 ( .A(n6187), .Y(n5996) );
  INVX3 U4036 ( .A(n5098), .Y(n5096) );
  CLKBUFX3 U4037 ( .A(n4302), .Y(n4298) );
  INVX12 U4038 ( .A(n5121), .Y(n5118) );
  CLKINVX1 U4039 ( .A(n8058), .Y(n8043) );
  NAND2X1 U4040 ( .A(n3410), .B(n6807), .Y(n8417) );
  OR2X1 U4041 ( .A(n6806), .B(n5475), .Y(n3410) );
  NAND2X1 U4042 ( .A(n3411), .B(n6810), .Y(n8418) );
  OR2X1 U4043 ( .A(n6809), .B(n5484), .Y(n3411) );
  AOI211X1 U4044 ( .A0(n5082), .A1(n5487), .B0(n6811), .C0(n6785), .Y(n6809)
         );
  NAND2X1 U4045 ( .A(n3412), .B(n6816), .Y(n8420) );
  OR2X1 U4046 ( .A(n6815), .B(n5502), .Y(n3412) );
  AOI211X1 U4047 ( .A0(n5082), .A1(n5505), .B0(n6817), .C0(n6785), .Y(n6815)
         );
  NAND2X1 U4048 ( .A(n3413), .B(n6873), .Y(n8439) );
  OR2X1 U4049 ( .A(n6872), .B(n5673), .Y(n3413) );
  AOI211X1 U4050 ( .A0(n5082), .A1(n5676), .B0(n6874), .C0(n6785), .Y(n6872)
         );
  NAND2X1 U4051 ( .A(n3414), .B(n6882), .Y(n8442) );
  OR2X1 U4052 ( .A(n6881), .B(n5700), .Y(n3414) );
  AOI211X1 U4053 ( .A0(n5082), .A1(n5703), .B0(n6883), .C0(n6785), .Y(n6881)
         );
  NAND2X1 U4054 ( .A(n3415), .B(n6888), .Y(n8444) );
  OR2X1 U4055 ( .A(n6887), .B(n5718), .Y(n3415) );
  AOI211X1 U4056 ( .A0(n5082), .A1(n5721), .B0(n6889), .C0(n6785), .Y(n6887)
         );
  NAND2X1 U4057 ( .A(n3416), .B(n6891), .Y(n8445) );
  OR2X1 U4058 ( .A(n6890), .B(n5727), .Y(n3416) );
  AOI211X1 U4059 ( .A0(n5082), .A1(n5730), .B0(n6892), .C0(n6785), .Y(n6890)
         );
  NAND2X1 U4060 ( .A(n3417), .B(n6837), .Y(n8427) );
  OR2X1 U4061 ( .A(n6836), .B(n5565), .Y(n3417) );
  AOI211X1 U4062 ( .A0(n5082), .A1(n5568), .B0(n6838), .C0(n6785), .Y(n6836)
         );
  NAND2X1 U4063 ( .A(n3418), .B(n6843), .Y(n8429) );
  OR2X1 U4064 ( .A(n6842), .B(n5583), .Y(n3418) );
  AOI211X1 U4065 ( .A0(n5082), .A1(n5586), .B0(n6844), .C0(n6785), .Y(n6842)
         );
  NAND2X1 U4066 ( .A(n3419), .B(n6846), .Y(n8430) );
  OR2X1 U4067 ( .A(n6845), .B(n5592), .Y(n3419) );
  AOI211X1 U4068 ( .A0(n5082), .A1(n5595), .B0(n6847), .C0(n6785), .Y(n6845)
         );
  NAND2X1 U4069 ( .A(n3420), .B(n6852), .Y(n8432) );
  OR2X1 U4070 ( .A(n6851), .B(n5610), .Y(n3420) );
  AOI211X1 U4071 ( .A0(n5082), .A1(n5613), .B0(n6853), .C0(n6785), .Y(n6851)
         );
  NAND2X1 U4072 ( .A(n3422), .B(n6825), .Y(n8423) );
  OR2X1 U4073 ( .A(n6824), .B(n5529), .Y(n3422) );
  AOI211X1 U4074 ( .A0(n5082), .A1(n5532), .B0(n6826), .C0(n6785), .Y(n6824)
         );
  NAND2X1 U4075 ( .A(n3423), .B(n6834), .Y(n8426) );
  OR2X1 U4076 ( .A(n6833), .B(n5556), .Y(n3423) );
  AOI211X1 U4077 ( .A0(n5082), .A1(n5559), .B0(n6835), .C0(n6785), .Y(n6833)
         );
  NAND2X1 U4078 ( .A(n3424), .B(n6840), .Y(n8428) );
  OR2X1 U4079 ( .A(n6839), .B(n5574), .Y(n3424) );
  AOI211X1 U4080 ( .A0(n5082), .A1(n5577), .B0(n6841), .C0(n6785), .Y(n6839)
         );
  NAND2X1 U4081 ( .A(n3425), .B(n6849), .Y(n8431) );
  OR2X1 U4082 ( .A(n6848), .B(n5601), .Y(n3425) );
  AOI211X1 U4083 ( .A0(n5082), .A1(n5604), .B0(n6850), .C0(n6785), .Y(n6848)
         );
  NAND2X1 U4084 ( .A(n3426), .B(n6855), .Y(n8433) );
  OR2X1 U4085 ( .A(n6854), .B(n5619), .Y(n3426) );
  AOI211X1 U4086 ( .A0(n5082), .A1(n5622), .B0(n6856), .C0(n6785), .Y(n6854)
         );
  NAND2X1 U4087 ( .A(n3430), .B(n6870), .Y(n8438) );
  OR2X1 U4088 ( .A(n6869), .B(n5664), .Y(n3430) );
  AOI211X1 U4089 ( .A0(n5082), .A1(n5667), .B0(n6871), .C0(n6785), .Y(n6869)
         );
  NAND2X1 U4090 ( .A(n3431), .B(n6879), .Y(n8441) );
  OR2X1 U4091 ( .A(n6878), .B(n5691), .Y(n3431) );
  AOI211X1 U4092 ( .A0(n5082), .A1(n5694), .B0(n6880), .C0(n6785), .Y(n6878)
         );
  NAND2X1 U4093 ( .A(n3432), .B(n6876), .Y(n8440) );
  OR2X1 U4094 ( .A(n6875), .B(n5682), .Y(n3432) );
  AOI211X1 U4095 ( .A0(n5082), .A1(n5685), .B0(n6877), .C0(n6785), .Y(n6875)
         );
  NAND2X1 U4096 ( .A(n3434), .B(n6885), .Y(n8443) );
  OR2X1 U4097 ( .A(n6884), .B(n5709), .Y(n3434) );
  AOI211X1 U4098 ( .A0(n5082), .A1(n5712), .B0(n6886), .C0(n6785), .Y(n6884)
         );
  NAND2X1 U4099 ( .A(n3468), .B(n5638), .Y(n8115) );
  OR2X1 U4100 ( .A(n5636), .B(n5637), .Y(n3468) );
  AOI211X1 U4101 ( .A0(n5100), .A1(n5640), .B0(n5641), .C0(n5414), .Y(n5636)
         );
  AOI211X1 U4102 ( .A0(n5072), .A1(n5892), .B0(n7885), .C0(n3357), .Y(n7880)
         );
  OAI21XL U4103 ( .A0(n7635), .A1(n5709), .B0(n7636), .Y(n8571) );
  AOI211X1 U4104 ( .A0(n5073), .A1(n5712), .B0(n7640), .C0(n7187), .Y(n7635)
         );
  AOI211X1 U4105 ( .A0(n5073), .A1(n5640), .B0(n7540), .C0(n7187), .Y(n7535)
         );
  NAND3X1 U4106 ( .A(n3462), .B(n3463), .C(n3464), .Y(n7337) );
  OAI21XL U4107 ( .A0(n6812), .A1(n5493), .B0(n6813), .Y(n8419) );
  OAI21XL U4108 ( .A0(n6974), .A1(n5979), .B0(n6975), .Y(n8473) );
  AOI211X1 U4109 ( .A0(n5072), .A1(n5874), .B0(n7863), .C0(n7187), .Y(n7858)
         );
  OAI222XL U4110 ( .A0(n5876), .A1(n5045), .B0(n5877), .B1(n5047), .C0(n5878), 
        .C1(n5050), .Y(n7863) );
  OAI21X1 U4111 ( .A0(n6938), .A1(n5871), .B0(n6939), .Y(n8461) );
  NOR2X1 U4112 ( .A(n3540), .B(n6785), .Y(n6938) );
  OAI21XL U4113 ( .A0(n7804), .A1(n5835), .B0(n7805), .Y(n8585) );
  AOI211X1 U4114 ( .A0(n5072), .A1(n5766), .B0(n7709), .C0(n7187), .Y(n7703)
         );
  OAI21X1 U4115 ( .A0(n6902), .A1(n5763), .B0(n6903), .Y(n8449) );
  NOR2X1 U4116 ( .A(n3539), .B(n6785), .Y(n6902) );
  OAI222XL U4117 ( .A0(n5732), .A1(n5045), .B0(n5733), .B1(n5047), .C0(n5734), 
        .C1(n5050), .Y(n7663) );
  OAI21XL U4118 ( .A0(n7603), .A1(n5691), .B0(n7604), .Y(n8569) );
  AOI211X1 U4119 ( .A0(n5073), .A1(n5694), .B0(n7608), .C0(n7187), .Y(n7603)
         );
  AOI211X1 U4120 ( .A0(n5073), .A1(n5658), .B0(n7563), .C0(n7187), .Y(n7558)
         );
  AOI211X1 U4121 ( .A0(n5073), .A1(n5622), .B0(n7507), .C0(n7187), .Y(n7500)
         );
  AOI211X1 U4122 ( .A0(n5073), .A1(n5586), .B0(n7460), .C0(n3357), .Y(n7455)
         );
  AOI211X1 U4123 ( .A0(n5073), .A1(n5514), .B0(n7360), .C0(n3358), .Y(n7355)
         );
  OAI21XL U4124 ( .A0(n6818), .A1(n5511), .B0(n6819), .Y(n8421) );
  AOI211X1 U4125 ( .A0(n5082), .A1(n5514), .B0(n6820), .C0(n6785), .Y(n6818)
         );
  AOI211X1 U4126 ( .A0(n5072), .A1(n5919), .B0(n7925), .C0(n3358), .Y(n7916)
         );
  OAI21XL U4127 ( .A0(n7669), .A1(n5736), .B0(n7670), .Y(n8574) );
  AOI211X1 U4128 ( .A0(n5072), .A1(n5739), .B0(n7674), .C0(n3357), .Y(n7669)
         );
  AOI211X1 U4129 ( .A0(n5073), .A1(n5595), .B0(n7471), .C0(n7187), .Y(n7466)
         );
  AOI211X1 U4130 ( .A0(n5074), .A1(n5451), .B0(n7258), .C0(n7187), .Y(n7251)
         );
  OAI222XL U4131 ( .A0(n5759), .A1(n5046), .B0(n5760), .B1(n5047), .C0(n5761), 
        .C1(n5050), .Y(n7697) );
  OAI222XL U4132 ( .A0(n5759), .A1(n5015), .B0(n5760), .B1(n5018), .C0(n5761), 
        .C1(n5023), .Y(n6901) );
  AOI211X1 U4133 ( .A0(n5073), .A1(n5685), .B0(n7597), .C0(n3357), .Y(n7592)
         );
  AOI211X1 U4134 ( .A0(n5073), .A1(n5613), .B0(n7494), .C0(n3358), .Y(n7489)
         );
  OAI222XL U4135 ( .A0(n5615), .A1(n5045), .B0(n5616), .B1(n5047), .C0(n5617), 
        .C1(n7189), .Y(n7494) );
  AOI211X1 U4136 ( .A0(n5073), .A1(n5541), .B0(n7394), .C0(n7187), .Y(n7389)
         );
  OAI21XL U4137 ( .A0(n7278), .A1(n5466), .B0(n7279), .Y(n8544) );
  OAI222XL U4138 ( .A0(n5966), .A1(n5029), .B0(n5967), .B1(n5031), .C0(n5968), 
        .C1(n5035), .Y(n7168) );
  OAI222XL U4139 ( .A0(n5966), .A1(n5004), .B0(n5967), .B1(n5005), .C0(n5968), 
        .C1(n5218), .Y(n6773) );
  OAI222XL U4140 ( .A0(n5966), .A1(n4990), .B0(n5967), .B1(n4992), .C0(n5968), 
        .C1(n4995), .Y(n6576) );
  OAI222XL U4141 ( .A0(n5966), .A1(n4979), .B0(n5967), .B1(n4980), .C0(n5968), 
        .C1(n4983), .Y(n6378) );
  OAI222XL U4142 ( .A0(n5966), .A1(n4963), .B0(n5967), .B1(n4967), .C0(n5968), 
        .C1(n4970), .Y(n6180) );
  OAI21X2 U4143 ( .A0(n5960), .A1(n5961), .B0(n5962), .Y(n8151) );
  AOI211X1 U4144 ( .A0(n5099), .A1(n5964), .B0(n5965), .C0(n5414), .Y(n5960)
         );
  OAI21X2 U4145 ( .A0(n5924), .A1(n5925), .B0(n5926), .Y(n8147) );
  AOI211X1 U4146 ( .A0(n5099), .A1(n5928), .B0(n5929), .C0(n5414), .Y(n5924)
         );
  AOI211X1 U4147 ( .A0(n5099), .A1(n5892), .B0(n5893), .C0(n5414), .Y(n5888)
         );
  AOI211X1 U4148 ( .A0(n5099), .A1(n5856), .B0(n5857), .C0(n5414), .Y(n5852)
         );
  AOI211X1 U4149 ( .A0(n5099), .A1(n5820), .B0(n5821), .C0(n5414), .Y(n5816)
         );
  AOI211X1 U4150 ( .A0(n5099), .A1(n5784), .B0(n5785), .C0(n5414), .Y(n5780)
         );
  AOI211X1 U4151 ( .A0(n5099), .A1(n5748), .B0(n5749), .C0(n5414), .Y(n5744)
         );
  AOI211X1 U4152 ( .A0(n5100), .A1(n5676), .B0(n5677), .C0(n5414), .Y(n5672)
         );
  NAND3X1 U4153 ( .A(n3453), .B(n3454), .C(n3455), .Y(n7012) );
  OAI21XL U4154 ( .A0(n6418), .A1(n5493), .B0(n6419), .Y(n8291) );
  NAND3X1 U4155 ( .A(n3450), .B(n3451), .C(n3452), .Y(n6222) );
  NAND3X1 U4156 ( .A(n3447), .B(n3448), .C(n3449), .Y(n6024) );
  AOI211X1 U4157 ( .A0(n5077), .A1(n5460), .B0(n7000), .C0(n6982), .Y(n6998)
         );
  OAI21XL U4158 ( .A0(n6406), .A1(n5457), .B0(n6407), .Y(n8287) );
  AOI211X1 U4159 ( .A0(n5101), .A1(n5460), .B0(n5461), .C0(n5414), .Y(n5456)
         );
  AOI211X1 U4160 ( .A0(n5077), .A1(n5424), .B0(n6988), .C0(n6982), .Y(n6986)
         );
  OAI21XL U4161 ( .A0(n6394), .A1(n5421), .B0(n6395), .Y(n8283) );
  AOI211X1 U4162 ( .A0(n5101), .A1(n5424), .B0(n5425), .C0(n5414), .Y(n5420)
         );
  OAI21XL U4163 ( .A0(n6184), .A1(n5979), .B0(n6185), .Y(n8217) );
  NOR2X1 U4164 ( .A(n3538), .B(n3364), .Y(n6184) );
  OAI21X2 U4165 ( .A0(n5942), .A1(n5943), .B0(n5944), .Y(n8149) );
  AOI211X1 U4166 ( .A0(n5099), .A1(n5946), .B0(n5947), .C0(n5414), .Y(n5942)
         );
  AOI211X1 U4167 ( .A0(n5099), .A1(n5910), .B0(n5911), .C0(n5414), .Y(n5906)
         );
  AOI211X1 U4168 ( .A0(n5099), .A1(n5838), .B0(n5839), .C0(n5414), .Y(n5834)
         );
  AOI211X1 U4169 ( .A0(n5099), .A1(n5766), .B0(n5767), .C0(n5414), .Y(n5762)
         );
  AOI211X1 U4170 ( .A0(n5100), .A1(n5730), .B0(n5731), .C0(n5414), .Y(n5726)
         );
  OAI21X2 U4171 ( .A0(n5654), .A1(n5655), .B0(n5656), .Y(n8117) );
  AOI211X1 U4172 ( .A0(n5100), .A1(n5658), .B0(n5659), .C0(n5414), .Y(n5654)
         );
  AOI211X1 U4173 ( .A0(n5100), .A1(n5586), .B0(n5587), .C0(n5414), .Y(n5582)
         );
  OAI21X2 U4174 ( .A0(n5546), .A1(n5547), .B0(n5548), .Y(n8105) );
  AOI211X1 U4175 ( .A0(n5100), .A1(n5550), .B0(n5551), .C0(n5414), .Y(n5546)
         );
  AOI211X1 U4176 ( .A0(n5076), .A1(n5514), .B0(n7018), .C0(n6982), .Y(n7016)
         );
  AOI211X1 U4177 ( .A0(n5100), .A1(n5514), .B0(n5515), .C0(n5414), .Y(n5510)
         );
  AOI211X1 U4178 ( .A0(n5100), .A1(n5478), .B0(n5479), .C0(n5414), .Y(n5474)
         );
  AOI211X1 U4179 ( .A0(n5077), .A1(n5442), .B0(n6994), .C0(n6982), .Y(n6992)
         );
  AOI211X1 U4180 ( .A0(n5101), .A1(n5442), .B0(n5443), .C0(n5414), .Y(n5438)
         );
  OAI21X2 U4181 ( .A0(n5951), .A1(n5952), .B0(n5953), .Y(n8150) );
  AOI211X1 U4182 ( .A0(n5099), .A1(n5955), .B0(n5956), .C0(n5414), .Y(n5951)
         );
  AOI211X1 U4183 ( .A0(n5099), .A1(n5919), .B0(n5920), .C0(n5414), .Y(n5915)
         );
  AOI211X1 U4184 ( .A0(n5099), .A1(n5883), .B0(n5884), .C0(n5414), .Y(n5879)
         );
  AOI211X1 U4185 ( .A0(n5099), .A1(n5847), .B0(n5848), .C0(n5414), .Y(n5843)
         );
  OAI21X2 U4186 ( .A0(n5807), .A1(n5808), .B0(n5809), .Y(n8134) );
  AOI211X1 U4187 ( .A0(n5099), .A1(n5811), .B0(n5812), .C0(n5414), .Y(n5807)
         );
  AOI211X1 U4188 ( .A0(n5099), .A1(n5775), .B0(n5776), .C0(n5414), .Y(n5771)
         );
  OAI21X2 U4189 ( .A0(n5735), .A1(n5736), .B0(n5737), .Y(n8126) );
  AOI211X1 U4190 ( .A0(n5099), .A1(n5739), .B0(n5740), .C0(n5414), .Y(n5735)
         );
  AOI211X1 U4191 ( .A0(n5100), .A1(n5703), .B0(n5704), .C0(n5414), .Y(n5699)
         );
  OAI21X2 U4192 ( .A0(n5663), .A1(n5664), .B0(n5665), .Y(n8118) );
  AOI211X1 U4193 ( .A0(n5100), .A1(n5667), .B0(n5668), .C0(n5414), .Y(n5663)
         );
  OAI21X2 U4194 ( .A0(n5627), .A1(n5628), .B0(n5629), .Y(n8114) );
  AOI211X1 U4195 ( .A0(n5100), .A1(n5631), .B0(n5632), .C0(n5414), .Y(n5627)
         );
  AOI211X1 U4196 ( .A0(n5100), .A1(n5595), .B0(n5596), .C0(n5414), .Y(n5591)
         );
  OAI21X2 U4197 ( .A0(n5555), .A1(n5556), .B0(n5557), .Y(n8106) );
  AOI211X1 U4198 ( .A0(n5100), .A1(n5559), .B0(n5560), .C0(n5414), .Y(n5555)
         );
  OAI21X2 U4199 ( .A0(n5519), .A1(n5520), .B0(n5521), .Y(n8102) );
  AOI211X1 U4200 ( .A0(n5100), .A1(n5523), .B0(n5524), .C0(n5414), .Y(n5519)
         );
  AOI211X1 U4201 ( .A0(n5100), .A1(n5487), .B0(n5488), .C0(n5414), .Y(n5483)
         );
  AOI211X1 U4202 ( .A0(n5077), .A1(n5451), .B0(n6997), .C0(n6982), .Y(n6995)
         );
  OAI21XL U4203 ( .A0(n6403), .A1(n5448), .B0(n6404), .Y(n8286) );
  AOI211X1 U4204 ( .A0(n5101), .A1(n5451), .B0(n5452), .C0(n5414), .Y(n5447)
         );
  OAI21XL U4205 ( .A0(n6386), .A1(n5408), .B0(n6387), .Y(n8282) );
  AOI211X1 U4206 ( .A0(n5091), .A1(n5412), .B0(n6389), .C0(n3356), .Y(n6386)
         );
  OAI21X2 U4207 ( .A0(n5407), .A1(n5408), .B0(n5409), .Y(n8090) );
  AOI211X1 U4208 ( .A0(n5101), .A1(n5412), .B0(n5413), .C0(n5414), .Y(n5407)
         );
  OAI21X2 U4209 ( .A0(n5969), .A1(n5970), .B0(n5971), .Y(n8152) );
  AOI211X1 U4210 ( .A0(n5099), .A1(n5973), .B0(n5974), .C0(n5414), .Y(n5969)
         );
  OAI21X2 U4211 ( .A0(n5933), .A1(n5934), .B0(n5935), .Y(n8148) );
  AOI211X1 U4212 ( .A0(n5099), .A1(n5937), .B0(n5938), .C0(n5414), .Y(n5933)
         );
  AOI211X1 U4213 ( .A0(n5099), .A1(n5901), .B0(n5902), .C0(n5414), .Y(n5897)
         );
  AOI211X1 U4214 ( .A0(n5099), .A1(n5865), .B0(n5866), .C0(n5414), .Y(n5861)
         );
  AOI211X1 U4215 ( .A0(n5099), .A1(n5829), .B0(n5830), .C0(n5414), .Y(n5825)
         );
  AOI211X1 U4216 ( .A0(n5099), .A1(n5793), .B0(n5794), .C0(n5414), .Y(n5789)
         );
  AOI211X1 U4217 ( .A0(n5099), .A1(n5757), .B0(n5758), .C0(n5414), .Y(n5753)
         );
  AOI211X1 U4218 ( .A0(n5100), .A1(n5721), .B0(n5722), .C0(n5414), .Y(n5717)
         );
  OAI21X2 U4219 ( .A0(n5681), .A1(n5682), .B0(n5683), .Y(n8120) );
  AOI211X1 U4220 ( .A0(n5100), .A1(n5685), .B0(n5686), .C0(n5414), .Y(n5681)
         );
  AOI211X1 U4221 ( .A0(n5100), .A1(n5649), .B0(n5650), .C0(n5414), .Y(n5645)
         );
  AOI211X1 U4222 ( .A0(n5100), .A1(n5613), .B0(n5614), .C0(n5414), .Y(n5609)
         );
  OAI21X2 U4223 ( .A0(n5573), .A1(n5574), .B0(n5575), .Y(n8108) );
  AOI211X1 U4224 ( .A0(n5100), .A1(n5577), .B0(n5578), .C0(n5414), .Y(n5573)
         );
  AOI211X1 U4225 ( .A0(n5076), .A1(n5541), .B0(n7027), .C0(n6982), .Y(n7025)
         );
  OAI21X2 U4226 ( .A0(n5537), .A1(n5538), .B0(n5539), .Y(n8104) );
  AOI211X1 U4227 ( .A0(n5100), .A1(n5541), .B0(n5542), .C0(n5414), .Y(n5537)
         );
  AOI211X1 U4228 ( .A0(n5100), .A1(n5505), .B0(n5506), .C0(n5414), .Y(n5501)
         );
  AOI211X1 U4229 ( .A0(n5077), .A1(n5469), .B0(n7003), .C0(n6982), .Y(n7001)
         );
  AOI211X1 U4230 ( .A0(n5101), .A1(n5469), .B0(n5470), .C0(n5414), .Y(n5465)
         );
  AOI211X1 U4231 ( .A0(n5077), .A1(n5433), .B0(n6991), .C0(n6982), .Y(n6989)
         );
  OAI21XL U4232 ( .A0(n6397), .A1(n5430), .B0(n6398), .Y(n8284) );
  AOI211X1 U4233 ( .A0(n5091), .A1(n5433), .B0(n6399), .C0(n3354), .Y(n6397)
         );
  AOI211X1 U4234 ( .A0(n5101), .A1(n5433), .B0(n5434), .C0(n5414), .Y(n5429)
         );
  INVX20 U4235 ( .A(n6977), .Y(n6785) );
  AND3X6 U4236 ( .A(n3542), .B(n3543), .C(n3544), .Y(n6977) );
  OAI33X1 U4237 ( .A0(n7191), .A1(n7192), .A2(n7184), .B0(n7193), .B1(n7194), 
        .B2(n5052), .Y(n7190) );
  OAI21X1 U4238 ( .A0(n5564), .A1(n5565), .B0(n5566), .Y(n8107) );
  OAI21X2 U4239 ( .A0(n5582), .A1(n5583), .B0(n5584), .Y(n8109) );
  OAI21X2 U4240 ( .A0(n5591), .A1(n5592), .B0(n5593), .Y(n8110) );
  OAI21X1 U4241 ( .A0(n6827), .A1(n5538), .B0(n6828), .Y(n8424) );
  OAI21X1 U4242 ( .A0(n6968), .A1(n5961), .B0(n6969), .Y(n8471) );
  OAI21X2 U4243 ( .A0(n5609), .A1(n5610), .B0(n5611), .Y(n8112) );
  OAI21X1 U4244 ( .A0(n6821), .A1(n5520), .B0(n6822), .Y(n8422) );
  OAI21X2 U4245 ( .A0(n5915), .A1(n5916), .B0(n5917), .Y(n8146) );
  OAI21X2 U4246 ( .A0(n5879), .A1(n5880), .B0(n5881), .Y(n8142) );
  OAI21X2 U4247 ( .A0(n5888), .A1(n5889), .B0(n5890), .Y(n8143) );
  OAI21X2 U4248 ( .A0(n5897), .A1(n5898), .B0(n5899), .Y(n8144) );
  OAI21X2 U4249 ( .A0(n5906), .A1(n5907), .B0(n5908), .Y(n8145) );
  INVX12 U4250 ( .A(n8020), .Y(n7187) );
  MX4X1 U4251 ( .A(n4047), .B(n4037), .C(n4042), .D(n4032), .S0(N2498), .S1(
        N2497), .Y(n3946) );
  CLKXOR2X8 U4252 ( .A(n4947), .B(\add_79/carry[5] ), .Y(N2498) );
  MX4XL U4253 ( .A(\ImageBuffer[0][3] ), .B(\ImageBuffer[1][3] ), .C(
        \ImageBuffer[2][3] ), .D(\ImageBuffer[3][3] ), .S0(n3486), .S1(n4306), 
        .Y(n4215) );
  MX4XL U4254 ( .A(\ImageBuffer[20][5] ), .B(\ImageBuffer[21][5] ), .C(
        \ImageBuffer[22][5] ), .D(\ImageBuffer[23][5] ), .S0(n3486), .S1(n3930), .Y(n3872) );
  MX4XL U4255 ( .A(\ImageBuffer[0][6] ), .B(\ImageBuffer[1][6] ), .C(
        \ImageBuffer[2][6] ), .D(\ImageBuffer[3][6] ), .S0(n3486), .S1(n3922), 
        .Y(n3898) );
  MX4XL U4256 ( .A(\ImageBuffer[56][6] ), .B(\ImageBuffer[57][6] ), .C(
        \ImageBuffer[58][6] ), .D(\ImageBuffer[59][6] ), .S0(n3486), .S1(n3922), .Y(n3881) );
  MX4XL U4257 ( .A(\ImageBuffer[48][6] ), .B(\ImageBuffer[49][6] ), .C(
        \ImageBuffer[50][6] ), .D(\ImageBuffer[51][6] ), .S0(n3935), .S1(n3920), .Y(n3883) );
  MX4XL U4258 ( .A(\ImageBuffer[52][6] ), .B(\ImageBuffer[53][6] ), .C(
        \ImageBuffer[54][6] ), .D(\ImageBuffer[55][6] ), .S0(n3940), .S1(n3923), .Y(n3882) );
  MX4XL U4259 ( .A(\ImageBuffer[44][6] ), .B(\ImageBuffer[45][6] ), .C(
        \ImageBuffer[46][6] ), .D(\ImageBuffer[47][6] ), .S0(n3935), .S1(n3929), .Y(n3885) );
  MX4X1 U4260 ( .A(\ImageBuffer[60][6] ), .B(\ImageBuffer[61][6] ), .C(
        \ImageBuffer[62][6] ), .D(\ImageBuffer[63][6] ), .S0(n3939), .S1(n3499), .Y(n3880) );
  BUFX4 U4261 ( .A(n3757), .Y(n3755) );
  CLKBUFX6 U4262 ( .A(n5123), .Y(n3920) );
  BUFX2 U4263 ( .A(n5119), .Y(n4302) );
  BUFX2 U4264 ( .A(n3366), .Y(n5059) );
  CLKINVX16 U4265 ( .A(n5124), .Y(n5123) );
  BUFX20 U4266 ( .A(n5123), .Y(n3932) );
  BUFX4 U4267 ( .A(n3924), .Y(n3925) );
  BUFX3 U4268 ( .A(n3923), .Y(n3928) );
  CLKINVX8 U4269 ( .A(n5126), .Y(n5125) );
  INVX3 U4270 ( .A(N2495), .Y(n5115) );
  BUFX4 U4271 ( .A(N2775), .Y(n4862) );
  BUFX4 U4272 ( .A(N2758), .Y(n4867) );
  BUFX8 U4273 ( .A(n3757), .Y(n3754) );
  BUFX12 U4274 ( .A(n4124), .Y(n4126) );
  AND2X2 U4275 ( .A(n8031), .B(n8029), .Y(n3366) );
  CLKBUFX2 U4276 ( .A(n5119), .Y(n3942) );
  BUFX16 U4277 ( .A(n4305), .Y(n4311) );
  CLKBUFX8 U4278 ( .A(n3932), .Y(n3921) );
  CLKBUFX2 U4279 ( .A(n3572), .Y(n5046) );
  BUFX12 U4280 ( .A(n4123), .Y(n4129) );
  BUFX6 U4281 ( .A(n3757), .Y(n4132) );
  CLKBUFX3 U4282 ( .A(n5121), .Y(n5119) );
  CLKBUFX2 U4283 ( .A(n4302), .Y(n4299) );
  BUFX8 U4284 ( .A(n4306), .Y(n4309) );
  BUFX8 U4285 ( .A(n4304), .Y(n4313) );
  INVX1 U4286 ( .A(n4864), .Y(n6393) );
  BUFX4 U4287 ( .A(n4317), .Y(n4308) );
  CLKBUFX8 U4288 ( .A(n4306), .Y(n4310) );
  INVX3 U4289 ( .A(N2488), .Y(n3479) );
  BUFX4 U4290 ( .A(N2495), .Y(n4135) );
  CLKBUFX8 U4291 ( .A(n5127), .Y(n3734) );
  CLKBUFX3 U4292 ( .A(n5064), .Y(n5062) );
  BUFX12 U4293 ( .A(n3936), .Y(n3938) );
  BUFX4 U4294 ( .A(n4303), .Y(n4314) );
  BUFX4 U4295 ( .A(n3924), .Y(n3926) );
  INVX1 U4296 ( .A(n4863), .Y(n6195) );
  INVXL U4297 ( .A(N2772), .Y(n6984) );
  INVXL U4298 ( .A(N2773), .Y(n7188) );
  INVX16 U4299 ( .A(n5128), .Y(n5127) );
  CLKBUFX3 U4300 ( .A(n5098), .Y(n5097) );
  INVX3 U4301 ( .A(N2490), .Y(n5122) );
  BUFX4 U4302 ( .A(n3757), .Y(n4128) );
  CLKBUFX3 U4303 ( .A(n5062), .Y(n5058) );
  INVX3 U4304 ( .A(N2489), .Y(n3408) );
  BUFX4 U4305 ( .A(n3922), .Y(n3930) );
  INVX3 U4306 ( .A(n3375), .Y(n3476) );
  OR2X2 U4307 ( .A(n4899), .B(n7196), .Y(n3367) );
  OR2X2 U4308 ( .A(n4926), .B(n7196), .Y(n3368) );
  OR2X2 U4309 ( .A(n7833), .B(n7196), .Y(n3369) );
  INVX12 U4310 ( .A(N2506), .Y(n3504) );
  BUFX8 U4311 ( .A(N2490), .Y(n3933) );
  NAND2X1 U4312 ( .A(n3443), .B(n5043), .Y(n7181) );
  BUFX6 U4313 ( .A(n5088), .Y(n5085) );
  MXI4X2 U4314 ( .A(n3553), .B(n3555), .C(n3554), .D(n3556), .S0(N2498), .S1(
        N2497), .Y(n3376) );
  BUFX4 U4315 ( .A(n3757), .Y(n4131) );
  BUFX4 U4316 ( .A(n3757), .Y(n3756) );
  BUFX4 U4317 ( .A(n3746), .Y(n3737) );
  OR3XL U4318 ( .A(n4311), .B(n4318), .C(n5118), .Y(n3370) );
  CLKBUFX3 U4319 ( .A(n5062), .Y(n5061) );
  CLKBUFX3 U4320 ( .A(n3923), .Y(n3499) );
  BUFX8 U4321 ( .A(n4305), .Y(n4312) );
  AND3X2 U4322 ( .A(n5126), .B(n7505), .C(n5128), .Y(n3371) );
  INVX3 U4323 ( .A(n3557), .Y(n7196) );
  OR2X1 U4324 ( .A(cmd[2]), .B(cmd[0]), .Y(n3372) );
  OR2X1 U4325 ( .A(cmd[2]), .B(cmd[1]), .Y(n3373) );
  INVX3 U4326 ( .A(n3550), .Y(n3944) );
  AND3X2 U4327 ( .A(n5405), .B(n5404), .C(cmd[3]), .Y(n3374) );
  NOR2BX1 U4328 ( .AN(n4863), .B(n4869), .Y(n5239) );
  OR3X2 U4329 ( .A(n5405), .B(cmd[2]), .C(n5404), .Y(n3375) );
  CLKINVX1 U4330 ( .A(n3570), .Y(N2505) );
  INVX3 U4331 ( .A(N2786), .Y(n5088) );
  MX4X1 U4332 ( .A(n3987), .B(n3977), .C(n3982), .D(n3972), .S0(N2498), .S1(
        N2497), .Y(n3943) );
  BUFX4 U4333 ( .A(n4134), .Y(n4122) );
  BUFX4 U4334 ( .A(n3748), .Y(n3750) );
  OAI221X1 U4335 ( .A0(n5115), .A1(n3348), .B0(n5112), .B1(n8063), .C0(n8069), 
        .Y(N2513) );
  BUFX4 U4336 ( .A(n4121), .Y(n4112) );
  OR3X2 U4337 ( .A(n5118), .B(n4318), .C(n3490), .Y(n3377) );
  OR3X2 U4338 ( .A(n5118), .B(n3409), .C(n3501), .Y(n3378) );
  OR3X2 U4339 ( .A(n3931), .B(n3409), .C(n5118), .Y(n3379) );
  OR3X2 U4340 ( .A(n3939), .B(n3409), .C(n3500), .Y(n3380) );
  OR3X2 U4341 ( .A(n3925), .B(n3409), .C(n3939), .Y(n3381) );
  BUFX4 U4342 ( .A(n5062), .Y(n5060) );
  OR3X2 U4343 ( .A(n5111), .B(n3491), .C(n3935), .Y(n3382) );
  BUFX8 U4344 ( .A(n3923), .Y(n3927) );
  CLKBUFX8 U4345 ( .A(n5093), .Y(n5092) );
  NAND3X1 U4346 ( .A(n3757), .B(n5118), .C(N2495), .Y(n3548) );
  NAND2X1 U4347 ( .A(n7967), .B(N2495), .Y(n3549) );
  CLKBUFX3 U4348 ( .A(n5113), .Y(n4307) );
  NAND3X1 U4349 ( .A(n5118), .B(n5117), .C(N2495), .Y(n3561) );
  NAND3X1 U4350 ( .A(n4300), .B(n5115), .C(n5116), .Y(n3562) );
  NAND3X1 U4351 ( .A(n5117), .B(n5115), .C(n5118), .Y(n3559) );
  NAND3X1 U4352 ( .A(n5117), .B(n5115), .C(n3939), .Y(n3558) );
  OR3X2 U4353 ( .A(n5118), .B(N2495), .C(n5117), .Y(n3383) );
  NAND2X1 U4354 ( .A(n8061), .B(n5400), .Y(n5982) );
  OAI32X4 U4355 ( .A0(n7595), .A1(n3352), .A2(n7596), .B0(n5060), .B1(n7602), 
        .Y(n5685) );
  OAI32X4 U4356 ( .A0(n7638), .A1(n3351), .A2(n7639), .B0(n5059), .B1(n7645), 
        .Y(n5712) );
  OAI32X1 U4357 ( .A0(n7971), .A1(n7192), .A2(n7965), .B0(n5067), .B1(n7928), 
        .Y(n7970) );
  CLKINVX1 U4358 ( .A(n7971), .Y(n7966) );
  NAND2X1 U4359 ( .A(n7934), .B(n7249), .Y(n7971) );
  INVX3 U4360 ( .A(n3380), .Y(n3391) );
  INVX3 U4361 ( .A(n3379), .Y(n3392) );
  INVX3 U4362 ( .A(n3370), .Y(n3393) );
  INVX3 U4363 ( .A(n3381), .Y(n3394) );
  INVX3 U4364 ( .A(n3378), .Y(n3395) );
  NOR3X2 U4365 ( .A(n7307), .B(N2490), .C(n7308), .Y(n7329) );
  INVX3 U4366 ( .A(N2491), .Y(n7307) );
  NOR3X2 U4367 ( .A(N2490), .B(N2491), .C(n7308), .Y(n7532) );
  INVX3 U4368 ( .A(N2492), .Y(n7308) );
  INVX3 U4369 ( .A(n3382), .Y(n3396) );
  INVX3 U4370 ( .A(n3377), .Y(n3397) );
  INVX3 U4371 ( .A(n3383), .Y(n3398) );
  NOR3X2 U4372 ( .A(n7310), .B(n5110), .C(n7311), .Y(n7204) );
  INVX3 U4373 ( .A(N2504), .Y(n7311) );
  INVX3 U4374 ( .A(N2503), .Y(n7310) );
  NOR3X2 U4375 ( .A(n5111), .B(n4310), .C(n3939), .Y(n7250) );
  INVX3 U4376 ( .A(n7395), .Y(n5545) );
  INVX3 U4377 ( .A(n7407), .Y(n5554) );
  INVX3 U4378 ( .A(n7438), .Y(n5572) );
  INVX3 U4379 ( .A(n7461), .Y(n5590) );
  INVX3 U4380 ( .A(n7472), .Y(n5599) );
  INVX3 U4381 ( .A(n7508), .Y(n5626) );
  INVX3 U4382 ( .A(n7541), .Y(n5644) );
  INVX3 U4383 ( .A(n7564), .Y(n5662) );
  INVX3 U4384 ( .A(n7575), .Y(n5671) );
  INVX3 U4385 ( .A(n7598), .Y(n5689) );
  OAI32X1 U4386 ( .A0(n7599), .A1(n7192), .A2(n7595), .B0(n3559), .B1(n7526), 
        .Y(n7598) );
  INVX3 U4387 ( .A(n7675), .Y(n5743) );
  OAI32X1 U4388 ( .A0(n7676), .A1(n7192), .A2(n7672), .B0(n3560), .B1(n4825), 
        .Y(n7675) );
  INVX3 U4389 ( .A(n7875), .Y(n5887) );
  NOR3X2 U4390 ( .A(N2503), .B(N2504), .C(n5110), .Y(n7834) );
  NOR3X2 U4391 ( .A(N2503), .B(N2504), .C(n5108), .Y(n7936) );
  AOI211XL U4392 ( .A0(n3398), .A1(n3371), .B0(n7990), .C0(n7991), .Y(n7989)
         );
  NOR3X2 U4393 ( .A(n3490), .B(n5118), .C(n5111), .Y(n7203) );
  NOR3X2 U4394 ( .A(n5118), .B(n4313), .C(n5111), .Y(n7235) );
  CLKBUFX3 U4395 ( .A(n5112), .Y(n5111) );
  NOR3X2 U4396 ( .A(n3939), .B(n4318), .C(n3491), .Y(n7277) );
  CLKBUFX3 U4397 ( .A(n3487), .Y(n4318) );
  NOR3X2 U4398 ( .A(n4309), .B(n4318), .C(n3939), .Y(n7309) );
  NAND2XL U4399 ( .A(n7331), .B(n3393), .Y(n7399) );
  NAND2XL U4400 ( .A(n7331), .B(n7250), .Y(n7365) );
  NOR3X2 U4401 ( .A(n7310), .B(n5108), .C(n7311), .Y(n7331) );
  NAND2XL U4402 ( .A(n7431), .B(n3393), .Y(n7499) );
  NAND2XL U4403 ( .A(n7431), .B(n3396), .Y(n7442) );
  NOR3X2 U4404 ( .A(n5109), .B(N2503), .C(n7311), .Y(n7431) );
  NAND2XL U4405 ( .A(n7534), .B(n3393), .Y(n7602) );
  NAND2XL U4406 ( .A(n7534), .B(n3397), .Y(n7579) );
  NOR3X2 U4407 ( .A(n5108), .B(N2503), .C(n7311), .Y(n7534) );
  NAND2XL U4408 ( .A(n7634), .B(n3397), .Y(n7679) );
  NAND2XL U4409 ( .A(n7634), .B(n3393), .Y(n7702) );
  NOR3X2 U4410 ( .A(n5109), .B(N2504), .C(n7310), .Y(n7634) );
  NAND2XL U4411 ( .A(n7735), .B(n3393), .Y(n7803) );
  NAND2XL U4412 ( .A(n7735), .B(n3396), .Y(n7746) );
  NOR3X2 U4413 ( .A(n5108), .B(N2504), .C(n7310), .Y(n7735) );
  NAND2X2 U4414 ( .A(n7179), .B(n4878), .Y(n5457) );
  NAND2X2 U4415 ( .A(n5041), .B(n4874), .Y(n5421) );
  NAND2X2 U4416 ( .A(n5044), .B(n4885), .Y(n5511) );
  NAND2X2 U4417 ( .A(n5043), .B(n4877), .Y(n5448) );
  NAND2X2 U4418 ( .A(n5044), .B(n4879), .Y(n5466) );
  NOR3X2 U4419 ( .A(n5118), .B(n3921), .C(n3408), .Y(n7234) );
  NOR3X2 U4420 ( .A(n3501), .B(n3939), .C(n3408), .Y(n7219) );
  NOR3X2 U4421 ( .A(n3939), .B(n3920), .C(n3408), .Y(n7249) );
  NOR3X2 U4422 ( .A(n7307), .B(n5122), .C(n7308), .Y(n7201) );
  NOR3X2 U4423 ( .A(n5122), .B(N2491), .C(n7308), .Y(n7429) );
  NOR3X2 U4424 ( .A(N2491), .B(N2492), .C(n5122), .Y(n7832) );
  NOR3X2 U4425 ( .A(n5122), .B(N2492), .C(n7307), .Y(n7632) );
  INVX12 U4434 ( .A(n3406), .Y(IRAM_D[7]) );
  NAND2X2 U4435 ( .A(n5043), .B(n4925), .Y(n5835) );
  NAND2X2 U4436 ( .A(n5044), .B(n4927), .Y(n5844) );
  NAND2X2 U4437 ( .A(n5044), .B(n4929), .Y(n5862) );
  NAND2X2 U4438 ( .A(n5044), .B(n4918), .Y(n5772) );
  NAND2X2 U4439 ( .A(n5044), .B(n4928), .Y(n5853) );
  NAND2X2 U4440 ( .A(n5044), .B(n4924), .Y(n5826) );
  NAND2X2 U4441 ( .A(n5044), .B(n4923), .Y(n5817) );
  NAND2X2 U4442 ( .A(n5044), .B(n4920), .Y(n5790) );
  NAND2X2 U4443 ( .A(n5044), .B(n4919), .Y(n5781) );
  NAND2X2 U4444 ( .A(n5044), .B(n4916), .Y(n5763) );
  INVX6 U4445 ( .A(n3408), .Y(n3409) );
  NAND2X2 U4446 ( .A(n5041), .B(n4880), .Y(n5475) );
  NAND2X2 U4447 ( .A(n7179), .B(n4882), .Y(n5484) );
  NAND2X2 U4448 ( .A(n7179), .B(n4884), .Y(n5502) );
  NAND2X2 U4449 ( .A(n5042), .B(n4905), .Y(n5673) );
  NAND2X2 U4450 ( .A(n5042), .B(n4909), .Y(n5700) );
  NAND2X2 U4451 ( .A(n5042), .B(n4911), .Y(n5718) );
  NAND2X2 U4452 ( .A(n5042), .B(n4912), .Y(n5727) );
  OR3X2 U4453 ( .A(n8018), .B(cmd[3]), .C(n8060), .Y(n3421) );
  NAND2X1 U4454 ( .A(n3421), .B(n8602), .Y(n8059) );
  NAND2X1 U4455 ( .A(N2748), .B(n4943), .Y(n3427) );
  NAND2X1 U4456 ( .A(sum[3]), .B(n5987), .Y(n3428) );
  NAND2X1 U4457 ( .A(N2756), .B(n5988), .Y(n3429) );
  AND3X2 U4458 ( .A(n3427), .B(n3428), .C(n3429), .Y(n7175) );
  NAND2X1 U4459 ( .A(n3433), .B(n5259), .Y(n5263) );
  OAI2BB1X1 U4460 ( .A0N(n5261), .A1N(n4873), .B0(n5077), .Y(n5260) );
  NAND3BX2 U4461 ( .AN(n5264), .B(n5263), .C(n5262), .Y(n5267) );
  AO21X1 U4462 ( .A0(n5082), .A1(n5541), .B0(n6829), .Y(n3435) );
  NOR2XL U4463 ( .A(n3435), .B(n6785), .Y(n6827) );
  AO21X1 U4464 ( .A0(n5082), .A1(n5523), .B0(n6823), .Y(n3436) );
  NOR2XL U4465 ( .A(n3436), .B(n6785), .Y(n6821) );
  AO21XL U4466 ( .A0(n5081), .A1(n5739), .B0(n6895), .Y(n3437) );
  NOR2XL U4467 ( .A(n3437), .B(n6785), .Y(n6893) );
  OAI32X4 U4468 ( .A0(n7672), .A1(n3352), .A2(n7673), .B0(n5059), .B1(n7679), 
        .Y(n5739) );
  AO21XL U4469 ( .A0(n5082), .A1(n5550), .B0(n6832), .Y(n3438) );
  NOR2XL U4470 ( .A(n3438), .B(n6785), .Y(n6830) );
  OAI32X4 U4471 ( .A0(n7403), .A1(n3351), .A2(n7404), .B0(n5061), .B1(n7412), 
        .Y(n5550) );
  AO21XL U4472 ( .A0(n5081), .A1(n5964), .B0(n6970), .Y(n3439) );
  NOR2XL U4473 ( .A(n3439), .B(n6785), .Y(n6968) );
  OAI32X4 U4474 ( .A0(n7990), .A1(n3351), .A2(n7991), .B0(n5061), .B1(n7997), 
        .Y(n5964) );
  OAI222XL U4475 ( .A0(n5966), .A1(n6786), .B0(n5967), .B1(n5019), .C0(n5968), 
        .C1(n5021), .Y(n6970) );
  NAND2X2 U4476 ( .A(N2749), .B(n4943), .Y(n3440) );
  NAND2X1 U4477 ( .A(sum[2]), .B(n5987), .Y(n3441) );
  MX4X1 U4478 ( .A(n4498), .B(n4488), .C(n4493), .D(n4483), .S0(N2516), .S1(
        N2515), .Y(N2757) );
  OR3X4 U4479 ( .A(n8013), .B(n3557), .C(n7304), .Y(n3443) );
  NAND2X1 U4480 ( .A(n3374), .B(n5406), .Y(n8031) );
  INVX4 U4481 ( .A(cmd[1]), .Y(n5405) );
  CLKINVX3 U4482 ( .A(cmd[2]), .Y(n5406) );
  NAND2X1 U4483 ( .A(N2746), .B(n4943), .Y(n3444) );
  NAND2X1 U4484 ( .A(sum[5]), .B(n5987), .Y(n3445) );
  NAND2X1 U4485 ( .A(N2754), .B(n5988), .Y(n3446) );
  BUFX4 U4486 ( .A(n5986), .Y(n4943) );
  NOR2X2 U4487 ( .A(n5405), .B(n3372), .Y(n8034) );
  BUFX4 U4488 ( .A(n8034), .Y(n3475) );
  NOR2X2 U4489 ( .A(n5404), .B(n3373), .Y(n8033) );
  BUFX4 U4490 ( .A(n8033), .Y(n3477) );
  OR2XL U4491 ( .A(n5498), .B(n4965), .Y(n3447) );
  OR2X1 U4492 ( .A(n5499), .B(n4969), .Y(n3448) );
  OR2X1 U4493 ( .A(n5500), .B(n4973), .Y(n3449) );
  OR2XL U4494 ( .A(n5498), .B(n4979), .Y(n3450) );
  OR2X1 U4495 ( .A(n5499), .B(n4981), .Y(n3451) );
  OR2X1 U4496 ( .A(n5500), .B(n4983), .Y(n3452) );
  OR2XL U4497 ( .A(n5498), .B(n6983), .Y(n3453) );
  OR2X1 U4498 ( .A(n5499), .B(n5034), .Y(n3454) );
  OR2X1 U4499 ( .A(n5500), .B(n5035), .Y(n3455) );
  OR2XL U4500 ( .A(n5498), .B(n5003), .Y(n3456) );
  OR2X1 U4501 ( .A(n5499), .B(n5006), .Y(n3457) );
  OR2X1 U4502 ( .A(n5500), .B(n5010), .Y(n3458) );
  NAND3X1 U4503 ( .A(n3456), .B(n3457), .C(n3458), .Y(n6617) );
  AO21XL U4504 ( .A0(n5074), .A1(n5424), .B0(n7213), .Y(n3459) );
  NOR2XL U4505 ( .A(n3459), .B(n7187), .Y(n7205) );
  OR2X2 U4506 ( .A(n7220), .B(n5430), .Y(n3460) );
  NAND2X2 U4507 ( .A(n3460), .B(n7221), .Y(n8540) );
  NAND2X2 U4508 ( .A(n5041), .B(n4875), .Y(n5430) );
  MXI2XL U4509 ( .A(\ImageBuffer[61][0] ), .B(n5040), .S0(n4875), .Y(n7221) );
  OR2X2 U4510 ( .A(n7236), .B(n5439), .Y(n3461) );
  NAND2X2 U4511 ( .A(n3461), .B(n7237), .Y(n8541) );
  NAND2X2 U4512 ( .A(n5042), .B(n4876), .Y(n5439) );
  MXI2XL U4513 ( .A(\ImageBuffer[60][0] ), .B(n5040), .S0(n4876), .Y(n7237) );
  OR2XL U4514 ( .A(n5498), .B(n5045), .Y(n3462) );
  OR2X1 U4515 ( .A(n5499), .B(n5048), .Y(n3463) );
  OR2XL U4516 ( .A(n5500), .B(n5049), .Y(n3464) );
  INVX3 U4517 ( .A(n7338), .Y(n5500) );
  AO21XL U4518 ( .A0(n5074), .A1(n5412), .B0(n7186), .Y(n3465) );
  NOR2XL U4519 ( .A(n3465), .B(n7187), .Y(n7176) );
  OAI222X1 U4520 ( .A0(n5415), .A1(n5045), .B0(n5416), .B1(n5047), .C0(n5418), 
        .C1(n5050), .Y(n7186) );
  AO21XL U4521 ( .A0(n5074), .A1(n5460), .B0(n7270), .Y(n3466) );
  NOR2X1 U4522 ( .A(n3466), .B(n3357), .Y(n7264) );
  OAI21XL U4523 ( .A0(n7264), .A1(n5457), .B0(n7265), .Y(n8543) );
  AO21XL U4524 ( .A0(n5074), .A1(n5469), .B0(n7285), .Y(n3467) );
  NOR2XL U4525 ( .A(n3467), .B(n7187), .Y(n7278) );
  BUFX20 U4526 ( .A(n3376), .Y(n5074) );
  MXI2XL U4527 ( .A(\ImageBuffer[38][7] ), .B(n4950), .S0(n4901), .Y(n5638) );
  AO21XL U4528 ( .A0(n5079), .A1(n5371), .B0(N2772), .Y(n5370) );
  NOR2BX1 U4529 ( .AN(N2773), .B(n5074), .Y(n5371) );
  MX4X2 U4530 ( .A(n4001), .B(n3999), .C(n4000), .D(n3998), .S0(n4108), .S1(
        n4135), .Y(n4002) );
  BUFX4 U4531 ( .A(n4110), .Y(n4108) );
  OAI32X1 U4532 ( .A0(n7807), .A1(n5057), .A2(n7808), .B0(n3351), .B1(n7815), 
        .Y(n7816) );
  NAND2X1 U4533 ( .A(n4865), .B(n6589), .Y(n5237) );
  BUFX4 U4534 ( .A(N2778), .Y(n4865) );
  OAI33X1 U4535 ( .A0(n7811), .A1(n7192), .A2(n7807), .B0(n3368), .B1(n7812), 
        .B2(n5071), .Y(n7810) );
  BUFX4 U4536 ( .A(n4297), .Y(n4301) );
  BUFX6 U4537 ( .A(n4299), .Y(n4300) );
  NOR2BX2 U4538 ( .AN(n4869), .B(n4863), .Y(n5147) );
  NOR2BX1 U4539 ( .AN(n4863), .B(n3361), .Y(n5332) );
  BUFX4 U4540 ( .A(N2776), .Y(n4863) );
  NOR4X1 U4541 ( .A(n5404), .B(n5406), .C(cmd[1]), .D(cmd[3]), .Y(n5986) );
  OAI211X2 U4542 ( .A0(n5232), .A1(n5155), .B0(n5129), .C0(n5138), .Y(n5130)
         );
  AND2X6 U4543 ( .A(n5131), .B(n5140), .Y(n5138) );
  NOR2BX1 U4544 ( .AN(n5091), .B(n4864), .Y(n5328) );
  BUFX4 U4545 ( .A(N2777), .Y(n4864) );
  AOI31X2 U4546 ( .A0(n5146), .A1(n5145), .A2(n5144), .B0(n5143), .Y(n5150) );
  NOR2X2 U4547 ( .A(n5132), .B(n5143), .Y(n5144) );
  BUFX12 U4548 ( .A(n7196), .Y(n5053) );
  AOI222X4 U4549 ( .A0(N2745), .A1(n4943), .B0(sum[6]), .B1(n5987), .C0(N2753), 
        .C1(n5988), .Y(n6583) );
  CLKBUFX3 U4550 ( .A(n5118), .Y(n3745) );
  INVX3 U4551 ( .A(n7909), .Y(n5914) );
  AOI211X2 U4552 ( .A0(n5195), .A1(n5207), .B0(n5194), .C0(n5210), .Y(n5196)
         );
  AOI31X4 U4553 ( .A0(n5209), .A1(n5208), .A2(n5207), .B0(n5206), .Y(n5213) );
  INVX3 U4554 ( .A(n7776), .Y(n5815) );
  AOI211X1 U4555 ( .A0(n5082), .A1(n5496), .B0(n6814), .C0(n6785), .Y(n6812)
         );
  AOI211XL U4556 ( .A0(n5090), .A1(n5496), .B0(n6420), .C0(n3355), .Y(n6418)
         );
  OAI32X4 U4557 ( .A0(n7335), .A1(n3352), .A2(n7336), .B0(n5061), .B1(n7342), 
        .Y(n5496) );
  NAND2X2 U4558 ( .A(N2770), .B(n5218), .Y(n5208) );
  NOR2X2 U4559 ( .A(n5218), .B(N2770), .Y(n5205) );
  INVX1 U4560 ( .A(n4865), .Y(n5218) );
  NAND2BX2 U4561 ( .AN(n5396), .B(n5378), .Y(n5391) );
  OAI31X4 U4562 ( .A0(n5397), .A1(n5396), .A2(n5395), .B0(n5394), .Y(N2708) );
  NOR2X1 U4563 ( .A(n5097), .B(N2767), .Y(n5396) );
  BUFX6 U4564 ( .A(\add_80/carry[2] ), .Y(n3470) );
  CLKINVX12 U4565 ( .A(n3504), .Y(n3474) );
  OAI221X4 U4566 ( .A0(n5117), .A1(n8076), .B0(n3491), .B1(n8077), .C0(n8084), 
        .Y(N2506) );
  MX4XL U4567 ( .A(\ImageBuffer[40][6] ), .B(\ImageBuffer[41][6] ), .C(
        \ImageBuffer[42][6] ), .D(\ImageBuffer[43][6] ), .S0(n4301), .S1(n4316), .Y(n4263) );
  MX4XL U4568 ( .A(\ImageBuffer[48][6] ), .B(\ImageBuffer[49][6] ), .C(
        \ImageBuffer[50][6] ), .D(\ImageBuffer[51][6] ), .S0(n4301), .S1(n4312), .Y(n4260) );
  MX4XL U4569 ( .A(\ImageBuffer[56][6] ), .B(\ImageBuffer[57][6] ), .C(
        \ImageBuffer[58][6] ), .D(\ImageBuffer[59][6] ), .S0(n4301), .S1(n5113), .Y(n4258) );
  MX4XL U4570 ( .A(\ImageBuffer[44][6] ), .B(\ImageBuffer[45][6] ), .C(
        \ImageBuffer[46][6] ), .D(\ImageBuffer[47][6] ), .S0(n4301), .S1(n4308), .Y(n4262) );
  MX4XL U4571 ( .A(\ImageBuffer[52][6] ), .B(\ImageBuffer[53][6] ), .C(
        \ImageBuffer[54][6] ), .D(\ImageBuffer[55][6] ), .S0(n4301), .S1(n4311), .Y(n4259) );
  MX4XL U4572 ( .A(\ImageBuffer[60][6] ), .B(\ImageBuffer[61][6] ), .C(
        \ImageBuffer[62][6] ), .D(\ImageBuffer[63][6] ), .S0(n4301), .S1(n4310), .Y(n4257) );
  NOR3BX4 U4573 ( .AN(n5270), .B(n5269), .C(n5255), .Y(n5256) );
  AOI211X2 U4574 ( .A0(n5254), .A1(n5265), .B0(n5357), .C0(n5268), .Y(n5255)
         );
  AOI31X2 U4575 ( .A0(n5189), .A1(n5166), .A2(n5182), .B0(n5185), .Y(n5167) );
  AOI211X2 U4576 ( .A0(n5133), .A1(n5144), .B0(n5132), .C0(n5147), .Y(n5134)
         );
  AOI31X2 U4577 ( .A0(n5145), .A1(n5131), .A2(n5130), .B0(n5142), .Y(n5133) );
  AO21XL U4578 ( .A0(n5079), .A1(n5342), .B0(n4873), .Y(n5341) );
  OAI211X1 U4579 ( .A0(n5342), .A1(n5079), .B0(n5341), .C0(n5351), .Y(n5343)
         );
  INVX20 U4580 ( .A(n5079), .Y(n5075) );
  AO21X2 U4581 ( .A0(n5079), .A1(n5313), .B0(n4866), .Y(n5312) );
  BUFX20 U4582 ( .A(n5080), .Y(n5079) );
  OAI21X2 U4583 ( .A0(n5429), .A1(n5430), .B0(n5431), .Y(n8092) );
  OAI21X2 U4584 ( .A0(n5834), .A1(n5835), .B0(n5836), .Y(n8137) );
  OAI21X2 U4585 ( .A0(n5510), .A1(n5511), .B0(n5512), .Y(n8101) );
  OAI21X2 U4586 ( .A0(n5726), .A1(n5727), .B0(n5728), .Y(n8125) );
  OAI21X2 U4587 ( .A0(n5753), .A1(n5754), .B0(n5755), .Y(n8128) );
  OAI21X2 U4588 ( .A0(n5762), .A1(n5763), .B0(n5764), .Y(n8129) );
  OAI21X4 U4589 ( .A0(n5600), .A1(n5601), .B0(n5602), .Y(n8111) );
  AOI211X4 U4590 ( .A0(n5100), .A1(n5604), .B0(n5605), .C0(n5414), .Y(n5600)
         );
  OAI21X4 U4591 ( .A0(n5690), .A1(n5691), .B0(n5692), .Y(n8121) );
  AOI211X4 U4592 ( .A0(n5100), .A1(n5694), .B0(n5695), .C0(n5414), .Y(n5690)
         );
  OAI21X2 U4593 ( .A0(n5717), .A1(n5718), .B0(n5719), .Y(n8124) );
  OAI21X2 U4594 ( .A0(n5744), .A1(n5745), .B0(n5746), .Y(n8127) );
  OAI21X2 U4595 ( .A0(n5780), .A1(n5781), .B0(n5782), .Y(n8131) );
  OAI21X2 U4596 ( .A0(n5789), .A1(n5790), .B0(n5791), .Y(n8132) );
  OAI21X4 U4597 ( .A0(n5798), .A1(n5799), .B0(n5800), .Y(n8133) );
  AOI211X4 U4598 ( .A0(n5099), .A1(n5802), .B0(n5803), .C0(n5414), .Y(n5798)
         );
  OAI21X2 U4599 ( .A0(n5816), .A1(n5817), .B0(n5818), .Y(n8135) );
  OAI21X2 U4600 ( .A0(n5825), .A1(n5826), .B0(n5827), .Y(n8136) );
  OAI21X2 U4601 ( .A0(n5852), .A1(n5853), .B0(n5854), .Y(n8139) );
  OAI21X4 U4602 ( .A0(n5870), .A1(n5871), .B0(n5872), .Y(n8141) );
  AOI211X4 U4603 ( .A0(n5099), .A1(n5874), .B0(n5875), .C0(n5414), .Y(n5870)
         );
  OAI21X2 U4604 ( .A0(n5483), .A1(n5484), .B0(n5485), .Y(n8098) );
  OAI21X2 U4605 ( .A0(n5699), .A1(n5700), .B0(n5701), .Y(n8122) );
  OAI21X2 U4606 ( .A0(n5771), .A1(n5772), .B0(n5773), .Y(n8130) );
  OAI21X2 U4607 ( .A0(n5501), .A1(n5502), .B0(n5503), .Y(n8100) );
  OAI21X2 U4608 ( .A0(n5474), .A1(n5475), .B0(n5476), .Y(n8097) );
  OAI21X4 U4609 ( .A0(n5528), .A1(n5529), .B0(n5530), .Y(n8103) );
  AOI211X4 U4610 ( .A0(n5100), .A1(n5532), .B0(n5533), .C0(n5414), .Y(n5528)
         );
  OAI21X2 U4611 ( .A0(n5456), .A1(n5457), .B0(n5458), .Y(n8095) );
  OAI21X4 U4612 ( .A0(n5618), .A1(n5619), .B0(n5620), .Y(n8113) );
  AOI211X4 U4613 ( .A0(n5100), .A1(n5622), .B0(n5623), .C0(n5414), .Y(n5618)
         );
  OAI21X2 U4614 ( .A0(n5861), .A1(n5862), .B0(n5863), .Y(n8140) );
  OAI21X2 U4615 ( .A0(n5843), .A1(n5844), .B0(n5845), .Y(n8138) );
  OAI21X2 U4616 ( .A0(n5438), .A1(n5439), .B0(n5440), .Y(n8093) );
  OAI21X2 U4617 ( .A0(n5420), .A1(n5421), .B0(n5422), .Y(n8091) );
  OAI21X2 U4618 ( .A0(n5447), .A1(n5448), .B0(n5449), .Y(n8094) );
  OAI21X2 U4619 ( .A0(n5465), .A1(n5466), .B0(n5467), .Y(n8096) );
  OAI21X2 U4620 ( .A0(n5645), .A1(n5646), .B0(n5647), .Y(n8116) );
  OAI21X2 U4621 ( .A0(n5672), .A1(n5673), .B0(n5674), .Y(n8119) );
  AOI31X2 U4622 ( .A0(n5267), .A1(n5266), .A2(n5265), .B0(n3492), .Y(n5271) );
  AOI31X2 U4623 ( .A0(n5266), .A1(n5253), .A2(n5252), .B0(n5264), .Y(n5254) );
  NAND2X1 U4624 ( .A(N2786), .B(n5277), .Y(n5266) );
  OR3X8 U4625 ( .A(n5167), .B(n5137), .C(n5199), .Y(n8088) );
  AOI31X4 U4626 ( .A0(n5158), .A1(n5136), .A2(n5151), .B0(n5154), .Y(n5137) );
  OAI21X4 U4627 ( .A0(n5492), .A1(n5493), .B0(n5494), .Y(n8099) );
  AOI211X4 U4628 ( .A0(n5100), .A1(n5496), .B0(n5497), .C0(n5414), .Y(n5492)
         );
  OAI21X4 U4629 ( .A0(n5708), .A1(n5709), .B0(n5710), .Y(n8123) );
  AOI211X4 U4630 ( .A0(n5100), .A1(n5712), .B0(n5713), .C0(n5414), .Y(n5708)
         );
  AO21X4 U4631 ( .A0(n5247), .A1(n5222), .B0(n4866), .Y(n5221) );
  AOI211X2 U4632 ( .A0(n5163), .A1(n5175), .B0(n5162), .C0(n5178), .Y(n5164)
         );
  AOI31X2 U4633 ( .A0(n5176), .A1(n5161), .A2(n5160), .B0(n5173), .Y(n5163) );
  BUFX12 U4634 ( .A(n8629), .Y(busy) );
  NOR2BX4 U4635 ( .AN(n5074), .B(N2781), .Y(n5324) );
  NOR3X2 U4636 ( .A(n5405), .B(cmd[3]), .C(n5406), .Y(n8021) );
  OAI222XL U4637 ( .A0(n5714), .A1(n5046), .B0(n5715), .B1(n5047), .C0(n5716), 
        .C1(n5050), .Y(n7640) );
  MX4X2 U4638 ( .A(n4532), .B(n4530), .C(n4531), .D(n4529), .S0(n3496), .S1(
        n4639), .Y(n4533) );
  MX4X2 U4639 ( .A(n4527), .B(n4525), .C(n4526), .D(n4524), .S0(n3496), .S1(
        n4639), .Y(n4528) );
  BUFX8 U4640 ( .A(n4641), .Y(n4639) );
  XNOR2X2 U4641 ( .A(\add_80/carry[3] ), .B(n5127), .Y(N2502) );
  XNOR2X2 U4642 ( .A(\add_80/carry[3] ), .B(n5127), .Y(n3493) );
  INVX8 U4643 ( .A(N2502), .Y(n5110) );
  BUFX20 U4644 ( .A(n5110), .Y(n5109) );
  OAI31X1 U4645 ( .A0(n5307), .A1(n5306), .A2(n5305), .B0(n5304), .Y(N2703) );
  NOR2X1 U4646 ( .A(n5310), .B(N2766), .Y(n5307) );
  INVX20 U4647 ( .A(n3545), .Y(n3505) );
  OAI21X4 U4648 ( .A0(n5120), .A1(n3348), .B0(n8071), .Y(n3545) );
  CLKINVX2 U4649 ( .A(n3479), .Y(n3480) );
  BUFX20 U4650 ( .A(n3941), .Y(n3486) );
  OR2X1 U4651 ( .A(n5127), .B(\add_80/carry[3] ), .Y(\add_80/carry[4] ) );
  AND2X6 U4652 ( .A(n3470), .B(N2495), .Y(\add_80/carry[3] ) );
  NAND2X1 U4653 ( .A(N2786), .B(n5186), .Y(n5176) );
  NOR2BX2 U4654 ( .AN(n5091), .B(n4870), .Y(n5357) );
  MX4XL U4655 ( .A(\ImageBuffer[28][4] ), .B(\ImageBuffer[29][4] ), .C(
        \ImageBuffer[30][4] ), .D(\ImageBuffer[31][4] ), .S0(n3742), .S1(n4125), .Y(n3663) );
  MX4XL U4656 ( .A(\ImageBuffer[20][4] ), .B(\ImageBuffer[21][4] ), .C(
        \ImageBuffer[22][4] ), .D(\ImageBuffer[23][4] ), .S0(n3742), .S1(n4130), .Y(n3665) );
  MX4XL U4657 ( .A(\ImageBuffer[36][4] ), .B(\ImageBuffer[37][4] ), .C(
        \ImageBuffer[38][4] ), .D(\ImageBuffer[39][4] ), .S0(n3742), .S1(n4125), .Y(n3660) );
  MX4XL U4658 ( .A(\ImageBuffer[24][4] ), .B(\ImageBuffer[25][4] ), .C(
        \ImageBuffer[26][4] ), .D(\ImageBuffer[27][4] ), .S0(n3742), .S1(n4129), .Y(n3664) );
  AOI211XL U4659 ( .A0(n5091), .A1(n5460), .B0(n6408), .C0(n3356), .Y(n6406)
         );
  AOI211XL U4660 ( .A0(n5091), .A1(n5442), .B0(n6402), .C0(n3354), .Y(n6400)
         );
  AOI211XL U4661 ( .A0(n5091), .A1(n5424), .B0(n6396), .C0(n3356), .Y(n6394)
         );
  AOI211XL U4662 ( .A0(n5091), .A1(n5469), .B0(n6411), .C0(n3354), .Y(n6409)
         );
  AOI211XL U4663 ( .A0(n5091), .A1(n5451), .B0(n6405), .C0(n3355), .Y(n6403)
         );
  NOR2BXL U4664 ( .AN(n4864), .B(n5091), .Y(n5316) );
  NOR2BXL U4665 ( .AN(N2769), .B(n5091), .Y(n5374) );
  NOR2BX1 U4666 ( .AN(n4864), .B(n5091), .Y(n5174) );
  NOR2BX1 U4667 ( .AN(n4870), .B(n5091), .Y(n5345) );
  NOR2BX4 U4668 ( .AN(N2765), .B(N2781), .Y(n5232) );
  BUFX8 U4669 ( .A(n3746), .Y(n3739) );
  CLKBUFX4 U4670 ( .A(n5128), .Y(n4109) );
  BUFX20 U4671 ( .A(n4118), .Y(n4117) );
  AOI2BB2XL U4672 ( .B0(n8079), .B1(n5127), .A0N(n5122), .A1N(n8080), .Y(n8082) );
  AOI2BB2XL U4673 ( .B0(n8065), .B1(n5127), .A0N(n5122), .A1N(n3523), .Y(n8068) );
  NOR2BX2 U4674 ( .AN(n5074), .B(N2765), .Y(n5353) );
  NAND2BX1 U4675 ( .AN(n4872), .B(n3944), .Y(n5253) );
  BUFX12 U4676 ( .A(N2763), .Y(n4872) );
  OAI21X1 U4677 ( .A0(n6893), .A1(n5736), .B0(n6894), .Y(n8446) );
  OAI21X1 U4678 ( .A0(n6830), .A1(n5547), .B0(n6831), .Y(n8425) );
  INVXL U4679 ( .A(n4308), .Y(n3490) );
  INVXL U4680 ( .A(n4305), .Y(n3491) );
  INVX16 U4681 ( .A(n5114), .Y(n5113) );
  BUFX20 U4682 ( .A(n5113), .Y(n4317) );
  BUFX16 U4683 ( .A(n4316), .Y(n4304) );
  BUFX20 U4684 ( .A(n4317), .Y(n4306) );
  BUFX20 U4685 ( .A(n4316), .Y(n4303) );
  BUFX16 U4686 ( .A(n4317), .Y(n4305) );
  BUFX4 U4687 ( .A(n4303), .Y(n4315) );
  BUFX4 U4688 ( .A(n3936), .Y(n3941) );
  BUFX16 U4689 ( .A(n3738), .Y(n3741) );
  MX4XL U4690 ( .A(\ImageBuffer[12][6] ), .B(\ImageBuffer[13][6] ), .C(
        \ImageBuffer[14][6] ), .D(\ImageBuffer[15][6] ), .S0(n4118), .S1(n4131), .Y(n4083) );
  MX4XL U4691 ( .A(\ImageBuffer[4][6] ), .B(\ImageBuffer[5][6] ), .C(
        \ImageBuffer[6][6] ), .D(\ImageBuffer[7][6] ), .S0(n4118), .S1(n4131), 
        .Y(n4085) );
  MX4X1 U4692 ( .A(\ImageBuffer[16][5] ), .B(\ImageBuffer[17][5] ), .C(
        \ImageBuffer[18][5] ), .D(\ImageBuffer[19][5] ), .S0(n3743), .S1(n3757), .Y(n3686) );
  NAND2BX4 U4693 ( .AN(n3361), .B(n4869), .Y(n5270) );
  NOR2BX4 U4694 ( .AN(N2768), .B(n5093), .Y(n5390) );
  NOR2BX4 U4695 ( .AN(n3361), .B(n4869), .Y(n5268) );
  NAND2BXL U4696 ( .AN(n3947), .B(n4863), .Y(n5180) );
  MX4X2 U4697 ( .A(n3778), .B(n3776), .C(n3777), .D(n3775), .S0(n3934), .S1(
        n3409), .Y(n3779) );
  NOR2BX4 U4698 ( .AN(n4870), .B(n4864), .Y(n5132) );
  NOR2BX2 U4699 ( .AN(n4864), .B(n4870), .Y(n5143) );
  AO21X2 U4700 ( .A0(n5155), .A1(n5232), .B0(n4873), .Y(n5129) );
  INVXL U4701 ( .A(n3487), .Y(n5112) );
  INVX16 U4702 ( .A(n7175), .Y(n6982) );
  INVX16 U4703 ( .A(n6780), .Y(n6588) );
  AOI211X1 U4704 ( .A0(n5092), .A1(n5983), .B0(n6384), .C0(n3350), .Y(n6382)
         );
  MX4XL U4705 ( .A(\ImageBuffer[52][0] ), .B(\ImageBuffer[53][0] ), .C(
        \ImageBuffer[54][0] ), .D(\ImageBuffer[55][0] ), .S0(n4114), .S1(n3747), .Y(n3952) );
  MX4X1 U4706 ( .A(n3606), .B(n3604), .C(n3605), .D(n3603), .S0(n3734), .S1(
        n3758), .Y(n3607) );
  MX4X2 U4707 ( .A(n3646), .B(n3644), .C(n3645), .D(n3643), .S0(n3734), .S1(
        n3758), .Y(n3647) );
  MX4X2 U4708 ( .A(n3641), .B(n3639), .C(n3640), .D(n3638), .S0(n3734), .S1(
        n3758), .Y(n3642) );
  CLKINVX20 U4709 ( .A(n5985), .Y(n5414) );
  AND3X8 U4710 ( .A(n3563), .B(n3564), .C(n3565), .Y(n5985) );
  AOI211X2 U4711 ( .A0(n5100), .A1(n5983), .B0(n5984), .C0(n5414), .Y(n5978)
         );
  INVXL U4712 ( .A(n3923), .Y(n3500) );
  INVXL U4713 ( .A(n3480), .Y(n3501) );
  CMPR22X2 U4714 ( .A(n3747), .B(n5118), .CO(\r2549/carry[2] ), .S(N2488) );
  BUFX20 U4715 ( .A(n3932), .Y(n3924) );
  CLKBUFX20 U4716 ( .A(n3932), .Y(n3923) );
  NAND2BX4 U4717 ( .AN(n8087), .B(n8086), .Y(n8076) );
  MXI2X2 U4718 ( .A(n8072), .B(n8065), .S0(n5118), .Y(n8071) );
  AOI2BB2X1 U4719 ( .B0(n8065), .B1(N2495), .A0N(n3408), .A1N(n3523), .Y(n8069) );
  INVX4 U4720 ( .A(n8075), .Y(n8065) );
  BUFX20 U4721 ( .A(n4112), .Y(n4115) );
  INVX3 U4722 ( .A(n3362), .Y(n3502) );
  AOI2BB1X4 U4723 ( .A0N(n5120), .A1N(n8076), .B0(n3571), .Y(n3570) );
  INVX6 U4724 ( .A(N2484), .Y(n5128) );
  CLKINVX16 U4725 ( .A(n3505), .Y(n3506) );
  BUFX20 U4726 ( .A(n3745), .Y(n3735) );
  CLKBUFX20 U4727 ( .A(n3739), .Y(n3740) );
  CLKBUFX4 U4728 ( .A(n5116), .Y(n3757) );
  CLKBUFX4 U4729 ( .A(n5116), .Y(n4134) );
  CLKBUFX4 U4730 ( .A(n5116), .Y(n3749) );
  BUFX12 U4731 ( .A(n4134), .Y(n4124) );
  BUFX20 U4732 ( .A(n4122), .Y(n4133) );
  BUFX20 U4733 ( .A(n3754), .Y(n4127) );
  CLKBUFX2 U4734 ( .A(n3747), .Y(n3752) );
  CLKBUFX2 U4735 ( .A(n3747), .Y(n3751) );
  BUFX12 U4736 ( .A(n3570), .Y(n3509) );
  BUFX6 U4737 ( .A(n3570), .Y(n3510) );
  CLKINVX12 U4738 ( .A(n3509), .Y(n3511) );
  CLKINVX12 U4739 ( .A(n3509), .Y(n3512) );
  CLKINVX12 U4740 ( .A(n3509), .Y(n3513) );
  CLKINVX12 U4741 ( .A(n3509), .Y(n3514) );
  CLKINVX8 U4742 ( .A(n3510), .Y(n3515) );
  CLKINVX8 U4743 ( .A(n3510), .Y(n3516) );
  CLKINVX8 U4744 ( .A(n3510), .Y(n3517) );
  CLKINVX8 U4745 ( .A(n3510), .Y(n3518) );
  CLKINVX8 U4746 ( .A(n3510), .Y(n3519) );
  BUFX8 U4747 ( .A(n8066), .Y(n3523) );
  AOI2BB2XL U4748 ( .B0(n8079), .B1(N2494), .A0N(n3500), .A1N(n8080), .Y(n8084) );
  NAND2X2 U4749 ( .A(n8080), .B(n8077), .Y(n8085) );
  AOI211X1 U4750 ( .A0(n5072), .A1(n5856), .B0(n7840), .C0(n3357), .Y(n7835)
         );
  OAI32X4 U4751 ( .A0(n7838), .A1(n3352), .A2(n7839), .B0(n5060), .B1(n7845), 
        .Y(n5856) );
  AOI211XL U4752 ( .A0(n5074), .A1(n5433), .B0(n7227), .C0(n3357), .Y(n7220)
         );
  OAI32X4 U4753 ( .A0(n7225), .A1(n3351), .A2(n7226), .B0(n5061), .B1(n7232), 
        .Y(n5433) );
  INVX8 U4754 ( .A(n7441), .Y(n5570) );
  OAI32X4 U4755 ( .A0(n7435), .A1(n5055), .A2(n7436), .B0(n3352), .B1(n7442), 
        .Y(n7441) );
  INVX8 U4756 ( .A(n7544), .Y(n5642) );
  OAI32X4 U4757 ( .A0(n7538), .A1(n5056), .A2(n7539), .B0(n3352), .B1(n7545), 
        .Y(n7544) );
  OAI32X4 U4758 ( .A0(n7358), .A1(n3351), .A2(n7359), .B0(n5061), .B1(n7365), 
        .Y(n5514) );
  OAI32X4 U4759 ( .A0(n7822), .A1(n3352), .A2(n7823), .B0(n5060), .B1(n7830), 
        .Y(n5847) );
  AOI211XL U4760 ( .A0(n5074), .A1(n5442), .B0(n7243), .C0(n3358), .Y(n7236)
         );
  OAI32X4 U4761 ( .A0(n7241), .A1(n3351), .A2(n7242), .B0(n5061), .B1(n7248), 
        .Y(n5442) );
  INVX3 U4762 ( .A(n8622), .Y(n7942) );
  OAI33X1 U4763 ( .A0(n7509), .A1(n5053), .A2(n7503), .B0(n7426), .B1(n7510), 
        .B2(n5071), .Y(n7512) );
  NAND2X2 U4764 ( .A(n7511), .B(n7304), .Y(n7426) );
  INVX8 U4765 ( .A(n7464), .Y(n5588) );
  OAI32X4 U4766 ( .A0(n7458), .A1(n5055), .A2(n7459), .B0(n3352), .B1(n7465), 
        .Y(n7464) );
  INVX8 U4767 ( .A(n7567), .Y(n5660) );
  OAI32X4 U4768 ( .A0(n7561), .A1(n5056), .A2(n7562), .B0(n3351), .B1(n7568), 
        .Y(n7567) );
  AOI211X1 U4769 ( .A0(n5072), .A1(n5757), .B0(n7697), .C0(n3357), .Y(n7692)
         );
  AOI211X1 U4770 ( .A0(n5081), .A1(n5757), .B0(n6901), .C0(n6785), .Y(n6899)
         );
  OAI32X4 U4771 ( .A0(n7695), .A1(n3351), .A2(n7696), .B0(n5060), .B1(n7702), 
        .Y(n5757) );
  OAI32X4 U4772 ( .A0(n7883), .A1(n3351), .A2(n7884), .B0(n5060), .B1(n7890), 
        .Y(n5892) );
  OAI32X4 U4773 ( .A0(n7906), .A1(n3351), .A2(n7907), .B0(n5055), .B1(n7914), 
        .Y(n5910) );
  OAI32X4 U4774 ( .A0(n7920), .A1(n3351), .A2(n7921), .B0(n5061), .B1(n7932), 
        .Y(n5919) );
  NAND3X2 U4775 ( .A(n7942), .B(n7954), .C(n7923), .Y(n7238) );
  NAND2X2 U4776 ( .A(n7980), .B(n7924), .Y(n7253) );
  OAI33X1 U4777 ( .A0(n7711), .A1(n7196), .A2(n7706), .B0(n7629), .B1(n7712), 
        .B2(n5071), .Y(n7714) );
  NAND2X2 U4778 ( .A(n7713), .B(n7304), .Y(n7629) );
  INVX8 U4779 ( .A(n7475), .Y(n5597) );
  OAI32X4 U4780 ( .A0(n7469), .A1(n5055), .A2(n7470), .B0(n3351), .B1(n7476), 
        .Y(n7475) );
  INVX8 U4781 ( .A(n7615), .Y(n5696) );
  OAI32X4 U4782 ( .A0(n7606), .A1(n5056), .A2(n7607), .B0(n3351), .B1(n7614), 
        .Y(n7615) );
  NOR2BX2 U4783 ( .AN(n7922), .B(n5115), .Y(n7182) );
  AOI211X1 U4784 ( .A0(n5073), .A1(n5730), .B0(n7663), .C0(n3358), .Y(n7658)
         );
  OAI32X4 U4785 ( .A0(n7661), .A1(n3352), .A2(n7662), .B0(n5059), .B1(n7668), 
        .Y(n5730) );
  AOI211X1 U4786 ( .A0(n5073), .A1(n5667), .B0(n7574), .C0(n7187), .Y(n7569)
         );
  OAI32X4 U4787 ( .A0(n7572), .A1(n3351), .A2(n7573), .B0(n5060), .B1(n7579), 
        .Y(n5667) );
  OAI32X4 U4788 ( .A0(n7392), .A1(n3352), .A2(n7393), .B0(n5061), .B1(n7399), 
        .Y(n5541) );
  OAI32X4 U4789 ( .A0(n7256), .A1(n3352), .A2(n7257), .B0(n5061), .B1(n7263), 
        .Y(n5451) );
  NAND3X2 U4790 ( .A(n7942), .B(n7954), .C(n7980), .Y(n7293) );
  INVX8 U4791 ( .A(n7413), .Y(n5552) );
  OAI32X4 U4792 ( .A0(n7403), .A1(n5055), .A2(n7404), .B0(n3352), .B1(n7412), 
        .Y(n7413) );
  INVX8 U4793 ( .A(n7578), .Y(n5669) );
  OAI32X4 U4794 ( .A0(n7572), .A1(n5056), .A2(n7573), .B0(n3352), .B1(n7579), 
        .Y(n7578) );
  INVX8 U4795 ( .A(n7779), .Y(n5813) );
  OAI32X4 U4796 ( .A0(n7773), .A1(n5057), .A2(n7774), .B0(n3352), .B1(n7780), 
        .Y(n7779) );
  OAI32X1 U4797 ( .A0(n7777), .A1(n7196), .A2(n7773), .B0(n3560), .B1(n7730), 
        .Y(n7778) );
  NAND2X2 U4798 ( .A(n7813), .B(n7304), .Y(n7730) );
  INVX3 U4799 ( .A(n7898), .Y(n5905) );
  OAI32XL U4800 ( .A0(n7899), .A1(n7192), .A2(n7895), .B0(n3559), .B1(n3369), 
        .Y(n7898) );
  BUFX12 U4801 ( .A(n8630), .Y(done) );
  MXI2X2 U4802 ( .A(reset), .B(n8039), .S0(n8038), .Y(n8037) );
  NOR2BX2 U4803 ( .AN(IRAM_valid), .B(reset), .Y(n8038) );
  NOR2BX2 U4804 ( .AN(n7967), .B(n5115), .Y(n7240) );
  OAI32X4 U4805 ( .A0(n7380), .A1(n3352), .A2(n7381), .B0(n5055), .B1(n7387), 
        .Y(n5532) );
  OAI33X1 U4806 ( .A0(n7384), .A1(n7192), .A2(n7380), .B0(n7323), .B1(n7385), 
        .B2(n5069), .Y(n7383) );
  OAI21X1 U4807 ( .A0(n5069), .A1(n4890), .B0(n7387), .Y(n7380) );
  OAI32X4 U4808 ( .A0(n7521), .A1(n3352), .A2(n7522), .B0(n5060), .B1(n7530), 
        .Y(n5631) );
  OAI21X1 U4809 ( .A0(n3548), .A1(n4908), .B0(n7530), .Y(n7521) );
  OAI32X4 U4810 ( .A0(n7446), .A1(n3351), .A2(n7447), .B0(n5060), .B1(n7453), 
        .Y(n5577) );
  OAI21X1 U4811 ( .A0(n5066), .A1(n4899), .B0(n7453), .Y(n7446) );
  AOI211X1 U4812 ( .A0(n5081), .A1(n5838), .B0(n6928), .C0(n6785), .Y(n6926)
         );
  AOI211X1 U4813 ( .A0(n5072), .A1(n5838), .B0(n7809), .C0(n3358), .Y(n7804)
         );
  OAI32X4 U4814 ( .A0(n7807), .A1(n3352), .A2(n7808), .B0(n5059), .B1(n7815), 
        .Y(n5838) );
  NOR3X2 U4815 ( .A(n3500), .B(n5118), .C(n3408), .Y(n7200) );
  OAI32X4 U4816 ( .A0(n7369), .A1(n3351), .A2(n7370), .B0(n5061), .B1(n7376), 
        .Y(n5523) );
  OAI32X4 U4817 ( .A0(n7503), .A1(n3351), .A2(n7504), .B0(n5060), .B1(n7513), 
        .Y(n5622) );
  OAI32X4 U4818 ( .A0(n7538), .A1(n3352), .A2(n7539), .B0(n5060), .B1(n7545), 
        .Y(n5640) );
  OAI32X4 U4819 ( .A0(n7268), .A1(n3352), .A2(n7269), .B0(n5061), .B1(n7275), 
        .Y(n5460) );
  NAND3X2 U4820 ( .A(n7506), .B(n7708), .C(n7405), .Y(n7918) );
  OAI33X4 U4821 ( .A0(n7553), .A1(n5053), .A2(n7549), .B0(n7529), .B1(n7554), 
        .B2(n5066), .Y(n7555) );
  OAI33X4 U4822 ( .A0(n7587), .A1(n5053), .A2(n7583), .B0(n7529), .B1(n7588), 
        .B2(n3562), .Y(n7589) );
  NAND2X2 U4823 ( .A(n7612), .B(n7304), .Y(n7529) );
  INVX8 U4824 ( .A(n7716), .Y(n5768) );
  OAI32X4 U4825 ( .A0(n7706), .A1(n5057), .A2(n7707), .B0(n3351), .B1(n7715), 
        .Y(n7716) );
  INVX8 U4826 ( .A(n7398), .Y(n5543) );
  OAI32X4 U4827 ( .A0(n7392), .A1(n5055), .A2(n7393), .B0(n3351), .B1(n7399), 
        .Y(n7398) );
  INVX8 U4828 ( .A(n7601), .Y(n5687) );
  OAI32X4 U4829 ( .A0(n7595), .A1(n5056), .A2(n7596), .B0(n3352), .B1(n7602), 
        .Y(n7601) );
  INVX3 U4830 ( .A(n7495), .Y(n5617) );
  BUFX12 U4831 ( .A(n8625), .Y(IRAM_A[3]) );
  OAI32X4 U4832 ( .A0(n7683), .A1(n3351), .A2(n7684), .B0(n5060), .B1(n7690), 
        .Y(n5748) );
  OAI21X1 U4833 ( .A0(n5069), .A1(n4917), .B0(n7690), .Y(n7683) );
  AOI211XL U4834 ( .A0(n7210), .A1(n3371), .B0(n7940), .C0(n7941), .Y(n7939)
         );
  OAI32X4 U4835 ( .A0(n7940), .A1(n3351), .A2(n7941), .B0(n5057), .B1(n7948), 
        .Y(n5928) );
  OAI32X1 U4836 ( .A0(n7945), .A1(n7192), .A2(n7940), .B0(n8057), .B1(n7928), 
        .Y(n7944) );
  OAI21X1 U4837 ( .A0(n5065), .A1(n7935), .B0(n7948), .Y(n7940) );
  AOI211XL U4838 ( .A0(n7418), .A1(n7182), .B0(n7419), .C0(n7420), .Y(n7417)
         );
  OAI32X4 U4839 ( .A0(n7419), .A1(n3351), .A2(n7420), .B0(n5056), .B1(n7427), 
        .Y(n5559) );
  OAI21X1 U4840 ( .A0(n5052), .A1(n4899), .B0(n7427), .Y(n7419) );
  OAI32X4 U4841 ( .A0(n7606), .A1(n3351), .A2(n7607), .B0(n5060), .B1(n7614), 
        .Y(n5694) );
  OAI32X4 U4842 ( .A0(n7952), .A1(n3352), .A2(n7953), .B0(n5059), .B1(n7960), 
        .Y(n5937) );
  OAI32X4 U4843 ( .A0(n7773), .A1(n3352), .A2(n7774), .B0(n5060), .B1(n7780), 
        .Y(n5811) );
  OAI32X4 U4844 ( .A0(n7283), .A1(n3352), .A2(n7284), .B0(n5061), .B1(n7290), 
        .Y(n5469) );
  AOI211XL U4845 ( .A0(n7224), .A1(n3371), .B0(n7952), .C0(n7953), .Y(n7951)
         );
  NOR3X2 U4846 ( .A(n3939), .B(n4125), .C(n5115), .Y(n7224) );
  NAND2XL U4847 ( .A(n7934), .B(n3391), .Y(n7994) );
  NAND2XL U4848 ( .A(n7934), .B(n7219), .Y(n7945) );
  NAND2XL U4849 ( .A(n7934), .B(n7234), .Y(n7957) );
  NAND2XL U4850 ( .A(n7934), .B(n3392), .Y(n8006) );
  NOR3X2 U4851 ( .A(N2491), .B(N2492), .C(N2490), .Y(n7934) );
  OAI33X1 U4852 ( .A0(n7910), .A1(n7196), .A2(n7906), .B0(n7829), .B1(n7911), 
        .B2(n5071), .Y(n7913) );
  OAI32X1 U4853 ( .A0(n7842), .A1(n7196), .A2(n7838), .B0(n5065), .B1(n7829), 
        .Y(n7843) );
  NAND2X2 U4854 ( .A(n7912), .B(n7304), .Y(n7829) );
  INVX3 U4855 ( .A(n7915), .Y(n5912) );
  INVX3 U4856 ( .A(n7998), .Y(n5966) );
  INVX8 U4857 ( .A(n7498), .Y(n5615) );
  OAI32X4 U4858 ( .A0(n7492), .A1(n5055), .A2(n7493), .B0(n3352), .B1(n7499), 
        .Y(n7498) );
  INVX8 U4859 ( .A(n7667), .Y(n5732) );
  OAI32X4 U4860 ( .A0(n7661), .A1(n5056), .A2(n7662), .B0(n3351), .B1(n7668), 
        .Y(n7667) );
  NAND2X2 U4861 ( .A(n7302), .B(n3557), .Y(n7193) );
  NAND2X4 U4862 ( .A(n8030), .B(n8031), .Y(n3557) );
  INVX3 U4863 ( .A(n7361), .Y(n5518) );
  INVX12 U4864 ( .A(n7708), .Y(IROM_A[5]) );
  INVX3 U4865 ( .A(n8617), .Y(n7708) );
  BUFX12 U4866 ( .A(n8627), .Y(IRAM_A[1]) );
  NOR2BX2 U4867 ( .AN(n7922), .B(N2495), .Y(n7255) );
  AOI211XL U4868 ( .A0(n3398), .A1(n7183), .B0(n7268), .C0(n7269), .Y(n7267)
         );
  AOI211XL U4869 ( .A0(n7224), .A1(n7183), .B0(n7225), .C0(n7226), .Y(n7223)
         );
  AOI211XL U4870 ( .A0(n7255), .A1(n7183), .B0(n7256), .C0(n7257), .Y(n7254)
         );
  NOR2X2 U4871 ( .A(n5128), .B(N2617), .Y(n7183) );
  OAI32X4 U4872 ( .A0(n7549), .A1(n3352), .A2(n7550), .B0(n5060), .B1(n7556), 
        .Y(n5649) );
  OAI21X1 U4873 ( .A0(n5066), .A1(n4908), .B0(n7556), .Y(n7549) );
  OAI32X4 U4874 ( .A0(n8002), .A1(n3352), .A2(n8003), .B0(n5061), .B1(n8009), 
        .Y(n5973) );
  OAI21X1 U4875 ( .A0(n5070), .A1(n7935), .B0(n8009), .Y(n8002) );
  OAI32X4 U4876 ( .A0(n7480), .A1(n3352), .A2(n7481), .B0(n5060), .B1(n7487), 
        .Y(n5604) );
  OAI21X1 U4877 ( .A0(n5069), .A1(n4899), .B0(n7487), .Y(n7480) );
  OAI32X4 U4878 ( .A0(n7723), .A1(n3352), .A2(n7724), .B0(n5059), .B1(n7731), 
        .Y(n5775) );
  OAI21X1 U4879 ( .A0(n5052), .A1(n4926), .B0(n7731), .Y(n7723) );
  OAI32X4 U4880 ( .A0(n7561), .A1(n3351), .A2(n7562), .B0(n5060), .B1(n7568), 
        .Y(n5658) );
  OAI32X4 U4881 ( .A0(n7796), .A1(n3351), .A2(n7797), .B0(n5060), .B1(n7803), 
        .Y(n5829) );
  OAI32X4 U4882 ( .A0(n7872), .A1(n3352), .A2(n7873), .B0(n5060), .B1(n7879), 
        .Y(n5883) );
  OAI32X4 U4883 ( .A0(n7458), .A1(n3352), .A2(n7459), .B0(n5061), .B1(n7465), 
        .Y(n5586) );
  OAI32X4 U4884 ( .A0(n7296), .A1(n3351), .A2(n7297), .B0(n5061), .B1(n7305), 
        .Y(n5478) );
  AOI211XL U4885 ( .A0(n7282), .A1(n3371), .B0(n8002), .C0(n8003), .Y(n8001)
         );
  AOI211XL U4886 ( .A0(n7282), .A1(n7183), .B0(n7283), .C0(n7284), .Y(n7281)
         );
  NOR3X2 U4887 ( .A(n4129), .B(N2495), .C(n3938), .Y(n7282) );
  AOI211X1 U4888 ( .A0(n7722), .A1(n7295), .B0(n7807), .C0(n7808), .Y(n7806)
         );
  AOI211XL U4889 ( .A0(n7722), .A1(n7255), .B0(n7773), .C0(n7774), .Y(n7772)
         );
  AOI211XL U4890 ( .A0(n7722), .A1(n7182), .B0(n7723), .C0(n7724), .Y(n7721)
         );
  AOI211XL U4891 ( .A0(n7722), .A1(n7282), .B0(n7796), .C0(n7797), .Y(n7795)
         );
  NOR3X2 U4892 ( .A(n5127), .B(n4947), .C(n5126), .Y(n7722) );
  AOI211XL U4893 ( .A0(n7418), .A1(n7240), .B0(n7458), .C0(n7459), .Y(n7457)
         );
  AOI211XL U4894 ( .A0(n7418), .A1(n7282), .B0(n7492), .C0(n7493), .Y(n7491)
         );
  AOI211XL U4895 ( .A0(n7418), .A1(n3398), .B0(n7480), .C0(n7481), .Y(n7479)
         );
  AOI211XL U4896 ( .A0(n7418), .A1(n7255), .B0(n7469), .C0(n7470), .Y(n7468)
         );
  NOR3X2 U4897 ( .A(n7505), .B(n5125), .C(n5128), .Y(n7418) );
  NAND2XL U4898 ( .A(n7733), .B(n3391), .Y(n7788) );
  NAND2XL U4899 ( .A(n7733), .B(n7234), .Y(n7754) );
  NAND2XL U4900 ( .A(n7733), .B(n3395), .Y(n7777) );
  NAND2XL U4901 ( .A(n7733), .B(n7200), .Y(n7727) );
  NAND2XL U4902 ( .A(n7733), .B(n3392), .Y(n7800) );
  NOR3X2 U4903 ( .A(N2490), .B(N2492), .C(n7307), .Y(n7733) );
  INVX3 U4904 ( .A(n7878), .Y(n5885) );
  INVX8 U4905 ( .A(n7514), .Y(n5624) );
  OAI32X4 U4906 ( .A0(n7503), .A1(n5055), .A2(n7504), .B0(n3351), .B1(n7513), 
        .Y(n7514) );
  INVX8 U4907 ( .A(n7678), .Y(n5741) );
  OAI32X4 U4908 ( .A0(n7672), .A1(n5056), .A2(n7673), .B0(n3351), .B1(n7679), 
        .Y(n7678) );
  NAND2X2 U4909 ( .A(n7302), .B(n7304), .Y(n7197) );
  INVX3 U4910 ( .A(n7372), .Y(n5527) );
  AOI211XL U4911 ( .A0(n7418), .A1(n7295), .B0(n7503), .C0(n7504), .Y(n7502)
         );
  AOI211XL U4912 ( .A0(n7183), .A1(n7295), .B0(n7296), .C0(n7297), .Y(n7294)
         );
  INVX3 U4913 ( .A(\sub_168_aco/B[0] ), .Y(n7295) );
  MXI2XL U4914 ( .A(n5401), .B(n5402), .S0(\state_cs[0] ), .Y(n5399) );
  NOR3X2 U4915 ( .A(n5401), .B(reset), .C(n4945), .Y(n8036) );
  NOR3BX1 U4916 ( .AN(n7924), .B(n7207), .C(n7968), .Y(n5401) );
  BUFX12 U4917 ( .A(n8628), .Y(IRAM_A[0]) );
  AOI211XL U4918 ( .A0(n7255), .A1(n3371), .B0(n7978), .C0(n7979), .Y(n7977)
         );
  OAI32X4 U4919 ( .A0(n7978), .A1(n3352), .A2(n7979), .B0(n5061), .B1(n7986), 
        .Y(n5955) );
  OAI21X1 U4920 ( .A0(n5068), .A1(n7935), .B0(n7986), .Y(n7978) );
  OAI32X4 U4921 ( .A0(n7583), .A1(n3351), .A2(n7584), .B0(n5060), .B1(n7590), 
        .Y(n5676) );
  OAI33X2 U4922 ( .A0(n7587), .A1(n7192), .A2(n7583), .B0(n7526), .B1(n7588), 
        .B2(n5069), .Y(n7586) );
  OAI21X1 U4923 ( .A0(n5069), .A1(n4908), .B0(n7590), .Y(n7583) );
  AOI211XL U4924 ( .A0(n7722), .A1(n7224), .B0(n7750), .C0(n7751), .Y(n7749)
         );
  OAI32X4 U4925 ( .A0(n7750), .A1(n3352), .A2(n7751), .B0(n5060), .B1(n7757), 
        .Y(n5793) );
  OAI21X1 U4926 ( .A0(n5066), .A1(n4926), .B0(n7757), .Y(n7750) );
  OAI32X4 U4927 ( .A0(n7621), .A1(n3352), .A2(n7622), .B0(n5059), .B1(n7630), 
        .Y(n5703) );
  OAI21X1 U4928 ( .A0(n5052), .A1(n4917), .B0(n7630), .Y(n7621) );
  OAI32X4 U4929 ( .A0(n7849), .A1(n3351), .A2(n7850), .B0(n5060), .B1(n7856), 
        .Y(n5865) );
  OAI32X4 U4930 ( .A0(n7435), .A1(n3352), .A2(n7436), .B0(n5061), .B1(n7442), 
        .Y(n5568) );
  OAI32X4 U4931 ( .A0(n7895), .A1(n3352), .A2(n7896), .B0(n5061), .B1(n7902), 
        .Y(n5901) );
  OAI32X4 U4932 ( .A0(n7469), .A1(n3351), .A2(n7470), .B0(n5060), .B1(n7476), 
        .Y(n5595) );
  OAI32X4 U4933 ( .A0(n7739), .A1(n3352), .A2(n7740), .B0(n5059), .B1(n7746), 
        .Y(n5784) );
  OAI32X4 U4934 ( .A0(n7346), .A1(n3351), .A2(n7347), .B0(n5061), .B1(n7353), 
        .Y(n5505) );
  OAI21X1 U4935 ( .A0(n5066), .A1(n4890), .B0(n7353), .Y(n7346) );
  INVX12 U4936 ( .A(n7954), .Y(IROM_A[1]) );
  NAND3X2 U4937 ( .A(n8621), .B(n7942), .C(n7923), .Y(n7208) );
  NAND3X2 U4938 ( .A(n8621), .B(n7942), .C(n7980), .Y(n7266) );
  INVX3 U4939 ( .A(n8621), .Y(n7954) );
  AOI211XL U4940 ( .A0(n7620), .A1(n3398), .B0(n7683), .C0(n7684), .Y(n7682)
         );
  AOI211XL U4941 ( .A0(n7620), .A1(n7182), .B0(n7621), .C0(n7622), .Y(n7619)
         );
  AOI211XL U4942 ( .A0(n7620), .A1(n7295), .B0(n7706), .C0(n7707), .Y(n7705)
         );
  AOI211XL U4943 ( .A0(n7620), .A1(n7282), .B0(n7695), .C0(n7696), .Y(n7694)
         );
  AOI211XL U4944 ( .A0(n7620), .A1(n7255), .B0(n7672), .C0(n7673), .Y(n7671)
         );
  NOR3X2 U4945 ( .A(n5126), .B(n4947), .C(n5128), .Y(n7620) );
  AOI211XL U4946 ( .A0(n7520), .A1(n7240), .B0(n7561), .C0(n7562), .Y(n7560)
         );
  AOI211XL U4947 ( .A0(n7520), .A1(n7295), .B0(n7606), .C0(n7607), .Y(n7605)
         );
  AOI211XL U4948 ( .A0(n7520), .A1(n3398), .B0(n7583), .C0(n7584), .Y(n7582)
         );
  AOI211XL U4949 ( .A0(n7520), .A1(n7224), .B0(n7549), .C0(n7550), .Y(n7548)
         );
  AOI211XL U4950 ( .A0(n7520), .A1(n7182), .B0(n7521), .C0(n7522), .Y(n7519)
         );
  NOR3X2 U4951 ( .A(n5127), .B(n5125), .C(n7505), .Y(n7520) );
  NAND2XL U4952 ( .A(n7832), .B(n3392), .Y(n7899) );
  NAND2XL U4953 ( .A(n7832), .B(n3395), .Y(n7876) );
  NAND2XL U4954 ( .A(n7832), .B(n7249), .Y(n7865) );
  NAND2XL U4955 ( .A(n7832), .B(n3394), .Y(n7910) );
  NAND2XL U4956 ( .A(n7832), .B(n7219), .Y(n7842) );
  NAND2XL U4957 ( .A(n7832), .B(n3391), .Y(n7887) );
  NAND3X2 U4958 ( .A(n7405), .B(n7506), .C(n8617), .Y(n7518) );
  OAI32X1 U4959 ( .A0(n7396), .A1(n5053), .A2(n7392), .B0(n3559), .B1(n7326), 
        .Y(n7397) );
  OAI32X1 U4960 ( .A0(n7373), .A1(n5053), .A2(n7369), .B0(n3560), .B1(n7326), 
        .Y(n7374) );
  OAI32X1 U4961 ( .A0(n7362), .A1(n5053), .A2(n7358), .B0(n3549), .B1(n7326), 
        .Y(n7363) );
  OAI32X1 U4962 ( .A0(n7339), .A1(n5053), .A2(n7335), .B0(n3547), .B1(n7326), 
        .Y(n7340) );
  NAND2X2 U4963 ( .A(n7410), .B(n7304), .Y(n7326) );
  INVX3 U4964 ( .A(n7901), .Y(n5903) );
  INVX8 U4965 ( .A(n7644), .Y(n5714) );
  OAI32X4 U4966 ( .A0(n7638), .A1(n5056), .A2(n7639), .B0(n3351), .B1(n7645), 
        .Y(n7644) );
  INVX8 U4967 ( .A(n7701), .Y(n5759) );
  OAI32X4 U4968 ( .A0(n7695), .A1(n5057), .A2(n7696), .B0(n3352), .B1(n7702), 
        .Y(n7701) );
  NAND2X2 U4969 ( .A(n8025), .B(n7304), .Y(n7931) );
  BUFX12 U4970 ( .A(n8624), .Y(IRAM_A[4]) );
  BUFX12 U4971 ( .A(n8626), .Y(IRAM_A[2]) );
  AND3XL U4972 ( .A(IRAM_A[1]), .B(IRAM_A[0]), .C(IRAM_A[2]), .Y(n8089) );
  BUFX12 U4973 ( .A(n8623), .Y(IRAM_A[5]) );
  AND4XL U4974 ( .A(IRAM_A[4]), .B(IRAM_A[3]), .C(IRAM_A[5]), .D(n8089), .Y(
        N13653) );
  AOI211XL U4975 ( .A0(n7317), .A1(n3398), .B0(n7380), .C0(n7381), .Y(n7379)
         );
  AOI211XL U4976 ( .A0(n7317), .A1(n7224), .B0(n7346), .C0(n7347), .Y(n7345)
         );
  AOI211XL U4977 ( .A0(n7317), .A1(n7182), .B0(n7318), .C0(n7319), .Y(n7316)
         );
  AOI211XL U4978 ( .A0(n7317), .A1(n7282), .B0(n7392), .C0(n7393), .Y(n7391)
         );
  AOI211XL U4979 ( .A0(n7317), .A1(n7240), .B0(n7358), .C0(n7359), .Y(n7357)
         );
  NOR2X2 U4980 ( .A(N2617), .B(n5127), .Y(n7317) );
  AOI211XL U4981 ( .A0(n7240), .A1(n3371), .B0(n7965), .C0(n7966), .Y(n7964)
         );
  OAI32X4 U4982 ( .A0(n7965), .A1(n3351), .A2(n7966), .B0(n5061), .B1(n7974), 
        .Y(n5946) );
  OAI21X1 U4983 ( .A0(n5067), .A1(n7935), .B0(n7974), .Y(n7965) );
  INVX12 U4984 ( .A(n7968), .Y(IROM_A[2]) );
  AOI211XL U4985 ( .A0(n7722), .A1(n3398), .B0(n7784), .C0(n7785), .Y(n7783)
         );
  OAI32X4 U4986 ( .A0(n7784), .A1(n3352), .A2(n7785), .B0(n5060), .B1(n7791), 
        .Y(n5820) );
  OAI21X1 U4987 ( .A0(n5069), .A1(n4926), .B0(n7791), .Y(n7784) );
  AOI211XL U4988 ( .A0(n7620), .A1(n7224), .B0(n7649), .C0(n7650), .Y(n7648)
         );
  OAI32X4 U4989 ( .A0(n7649), .A1(n3351), .A2(n7650), .B0(n5060), .B1(n7656), 
        .Y(n5721) );
  OAI21X1 U4990 ( .A0(n5066), .A1(n4917), .B0(n7656), .Y(n7649) );
  AOI211XL U4991 ( .A0(n7182), .A1(n7183), .B0(n7184), .C0(n7185), .Y(n7180)
         );
  OAI32X4 U4992 ( .A0(n7184), .A1(n3351), .A2(n7185), .B0(n5060), .B1(n7198), 
        .Y(n5412) );
  OAI21X1 U4993 ( .A0(n4881), .A1(n5052), .B0(n7198), .Y(n7184) );
  OAI32X4 U4994 ( .A0(n7492), .A1(n3351), .A2(n7493), .B0(n5060), .B1(n7499), 
        .Y(n5613) );
  OAI32X4 U4995 ( .A0(n7211), .A1(n3352), .A2(n7212), .B0(n5060), .B1(n7218), 
        .Y(n5424) );
  OAI32X4 U4996 ( .A0(n7318), .A1(n3351), .A2(n7319), .B0(n5061), .B1(n7327), 
        .Y(n5487) );
  OAI21X1 U4997 ( .A0(n5052), .A1(n4890), .B0(n7327), .Y(n7318) );
  OAI32X4 U4998 ( .A0(n7762), .A1(n3351), .A2(n7763), .B0(n5059), .B1(n7769), 
        .Y(n5802) );
  AOI211XL U4999 ( .A0(n7821), .A1(n7295), .B0(n7906), .C0(n7907), .Y(n7905)
         );
  AOI211XL U5000 ( .A0(n7821), .A1(n3398), .B0(n7883), .C0(n7884), .Y(n7882)
         );
  AOI211XL U5001 ( .A0(n7821), .A1(n7282), .B0(n7895), .C0(n7896), .Y(n7894)
         );
  AOI211XL U5002 ( .A0(n7821), .A1(n7255), .B0(n7872), .C0(n7873), .Y(n7871)
         );
  AOI211XL U5003 ( .A0(n7821), .A1(n7240), .B0(n7861), .C0(n7862), .Y(n7860)
         );
  AOI211XL U5004 ( .A0(n7821), .A1(n7224), .B0(n7849), .C0(n7850), .Y(n7848)
         );
  NOR3X2 U5005 ( .A(n5125), .B(n4947), .C(n5128), .Y(n7821) );
  INVX12 U5006 ( .A(n7942), .Y(IROM_A[0]) );
  NAND3X2 U5007 ( .A(n8622), .B(n7954), .C(n7923), .Y(n7222) );
  NAND3X2 U5008 ( .A(n8622), .B(n7954), .C(n7980), .Y(n7280) );
  INVX12 U5009 ( .A(n7506), .Y(IROM_A[4]) );
  NAND3X2 U5010 ( .A(n8618), .B(n7405), .C(n8617), .Y(n7314) );
  NAND3X2 U5011 ( .A(n7405), .B(n7708), .C(n8618), .Y(n7720) );
  INVX3 U5012 ( .A(n8618), .Y(n7506) );
  INVX12 U5013 ( .A(n7405), .Y(IROM_A[3]) );
  NAND3X2 U5014 ( .A(n8619), .B(n7506), .C(n8617), .Y(n7416) );
  NAND3X2 U5015 ( .A(n8619), .B(n7708), .C(n8618), .Y(n7618) );
  NAND3X2 U5016 ( .A(n7506), .B(n7708), .C(n8619), .Y(n7819) );
  NAND3X2 U5017 ( .A(n8618), .B(n8619), .C(n8617), .Y(n7207) );
  INVX3 U5018 ( .A(n8619), .Y(n7405) );
  NAND2XL U5019 ( .A(n7632), .B(n7219), .Y(n7642) );
  NAND2XL U5020 ( .A(n7632), .B(n3392), .Y(n7699) );
  NAND2XL U5021 ( .A(n7632), .B(n3395), .Y(n7676) );
  NAND2XL U5022 ( .A(n7632), .B(n7249), .Y(n7665) );
  NAND2XL U5023 ( .A(n7632), .B(n3394), .Y(n7711) );
  NAND2XL U5024 ( .A(n7632), .B(n3391), .Y(n7687) );
  AO21XL U5025 ( .A0(n5095), .A1(n5983), .B0(n6186), .Y(n3538) );
  OAI32X4 U5026 ( .A0(n8016), .A1(n3351), .A2(n8017), .B0(n5058), .B1(n8027), 
        .Y(n5983) );
  AO21XL U5027 ( .A0(n5081), .A1(n5766), .B0(n6904), .Y(n3539) );
  OAI32X4 U5028 ( .A0(n7706), .A1(n3352), .A2(n7707), .B0(n5059), .B1(n7715), 
        .Y(n5766) );
  AO21XL U5029 ( .A0(n5081), .A1(n5874), .B0(n6940), .Y(n3540) );
  OAI32X4 U5030 ( .A0(n7861), .A1(n3352), .A2(n7862), .B0(n5060), .B1(n7868), 
        .Y(n5874) );
  INVX1 U5031 ( .A(n7524), .Y(n5635) );
  CLKBUFX2 U5032 ( .A(n3746), .Y(n3738) );
  INVX3 U5033 ( .A(n7483), .Y(n5608) );
  INVX3 U5034 ( .A(n7383), .Y(n5536) );
  INVX1 U5035 ( .A(n8007), .Y(n5976) );
  INVX1 U5036 ( .A(n7984), .Y(n5958) );
  INVX1 U5037 ( .A(n7972), .Y(n5949) );
  INVX1 U5038 ( .A(n7946), .Y(n5931) );
  INVX1 U5039 ( .A(n7586), .Y(n5680) );
  INVX1 U5040 ( .A(n7552), .Y(n5653) );
  CLKBUFX3 U5041 ( .A(n5062), .Y(n5057) );
  BUFX4 U5042 ( .A(N2495), .Y(n3758) );
  OAI33X1 U5043 ( .A0(n7610), .A1(n7192), .A2(n7606), .B0(n7526), .B1(n7611), 
        .B2(n5071), .Y(n7609) );
  NOR2BX1 U5044 ( .AN(n3947), .B(n4863), .Y(n5178) );
  NAND2X1 U5045 ( .A(N2767), .B(n5219), .Y(n5198) );
  NAND2BX1 U5046 ( .AN(N2779), .B(n3944), .Y(n5161) );
  INVX12 U5047 ( .A(n3551), .Y(N2781) );
  MX4XL U5048 ( .A(\ImageBuffer[12][1] ), .B(\ImageBuffer[13][1] ), .C(
        \ImageBuffer[14][1] ), .D(\ImageBuffer[15][1] ), .S0(n5120), .S1(n3920), .Y(n3795) );
  MX4XL U5049 ( .A(\ImageBuffer[44][1] ), .B(\ImageBuffer[45][1] ), .C(
        \ImageBuffer[46][1] ), .D(\ImageBuffer[47][1] ), .S0(n3939), .S1(n3925), .Y(n3785) );
  MX4XL U5050 ( .A(\ImageBuffer[48][7] ), .B(\ImageBuffer[49][7] ), .C(
        \ImageBuffer[50][7] ), .D(\ImageBuffer[51][7] ), .S0(n3938), .S1(n3932), .Y(n3903) );
  NOR2BX2 U5051 ( .AN(N2768), .B(n4863), .Y(n5210) );
  INVX1 U5052 ( .A(n7930), .Y(n5922) );
  INVX1 U5053 ( .A(n7855), .Y(n5868) );
  NAND2BXL U5054 ( .AN(n5277), .B(n5085), .Y(n3541) );
  MX4X1 U5055 ( .A(n3823), .B(n3821), .C(n3822), .D(n3820), .S0(n3933), .S1(
        n3409), .Y(n3824) );
  MX4XL U5056 ( .A(\ImageBuffer[28][1] ), .B(\ImageBuffer[29][1] ), .C(
        \ImageBuffer[30][1] ), .D(\ImageBuffer[31][1] ), .S0(n4115), .S1(n4126), .Y(n3978) );
  MX4XL U5057 ( .A(\ImageBuffer[40][2] ), .B(\ImageBuffer[41][2] ), .C(
        \ImageBuffer[42][2] ), .D(\ImageBuffer[43][2] ), .S0(n3506), .S1(n3485), .Y(n4525) );
  MX4XL U5058 ( .A(\ImageBuffer[56][3] ), .B(\ImageBuffer[57][3] ), .C(
        \ImageBuffer[58][3] ), .D(\ImageBuffer[59][3] ), .S0(n3347), .S1(n3483), .Y(n4540) );
  MX4XL U5059 ( .A(\ImageBuffer[16][2] ), .B(\ImageBuffer[17][2] ), .C(
        \ImageBuffer[18][2] ), .D(\ImageBuffer[19][2] ), .S0(n3342), .S1(n3482), .Y(n4532) );
  MX4XL U5060 ( .A(\ImageBuffer[32][2] ), .B(\ImageBuffer[33][2] ), .C(
        \ImageBuffer[34][2] ), .D(\ImageBuffer[35][2] ), .S0(n3342), .S1(n3482), .Y(n4527) );
  MX4XL U5061 ( .A(\ImageBuffer[36][2] ), .B(\ImageBuffer[37][2] ), .C(
        \ImageBuffer[38][2] ), .D(\ImageBuffer[39][2] ), .S0(n3346), .S1(n3484), .Y(n4526) );
  CLKBUFX2 U5062 ( .A(n4121), .Y(n4113) );
  INVX3 U5063 ( .A(n5289), .Y(N2675) );
  NOR2BX1 U5064 ( .AN(N2765), .B(n5074), .Y(n5261) );
  CLKMX2X6 U5065 ( .A(n8085), .B(n8079), .S0(n5118), .Y(n3571) );
  NOR2BX1 U5066 ( .AN(n5118), .B(n5117), .Y(\add_80/carry[2] ) );
  MX4XL U5067 ( .A(\ImageBuffer[4][5] ), .B(\ImageBuffer[5][5] ), .C(
        \ImageBuffer[6][5] ), .D(\ImageBuffer[7][5] ), .S0(n4300), .S1(n3926), 
        .Y(n3877) );
  MX4XL U5068 ( .A(\ImageBuffer[12][5] ), .B(\ImageBuffer[13][5] ), .C(
        \ImageBuffer[14][5] ), .D(\ImageBuffer[15][5] ), .S0(n4300), .S1(n3924), .Y(n3875) );
  INVX4 U5069 ( .A(n7388), .Y(n5534) );
  INVX1 U5070 ( .A(n7982), .Y(n5959) );
  INVX1 U5071 ( .A(n7970), .Y(n5950) );
  INVX1 U5072 ( .A(n7944), .Y(n5932) );
  INVX1 U5073 ( .A(n7286), .Y(n5473) );
  INVX1 U5074 ( .A(n7259), .Y(n5455) );
  INVX1 U5075 ( .A(n7244), .Y(n5446) );
  INVX1 U5076 ( .A(n7214), .Y(n5428) );
  INVX1 U5077 ( .A(n7288), .Y(n5472) );
  INVX1 U5078 ( .A(n7261), .Y(n5454) );
  INVX1 U5079 ( .A(n7246), .Y(n5445) );
  INVX1 U5080 ( .A(n7216), .Y(n5427) );
  OAI31X2 U5081 ( .A0(n5339), .A1(n5338), .A2(n5337), .B0(n5336), .Y(N2706) );
  NOR2X2 U5082 ( .A(n5186), .B(N2786), .Y(n5173) );
  NOR2X2 U5083 ( .A(n5187), .B(n4868), .Y(n5153) );
  NOR2X1 U5084 ( .A(n5188), .B(N2766), .Y(n5217) );
  NOR2BX1 U5085 ( .AN(N2781), .B(n5074), .Y(n5170) );
  NAND2X2 U5086 ( .A(N2755), .B(n5988), .Y(n3544) );
  CLKINVX4 U5087 ( .A(n3967), .Y(n3553) );
  AND2X2 U5088 ( .A(\add_80/carry[4] ), .B(n5125), .Y(\add_80/carry[5] ) );
  INVX12 U5089 ( .A(n3552), .Y(N2779) );
  CLKINVX8 U5090 ( .A(n3943), .Y(n5080) );
  MX4X4 U5091 ( .A(n3986), .B(n3984), .C(n3985), .D(n3983), .S0(n4108), .S1(
        n4135), .Y(n3987) );
  MX4XL U5092 ( .A(\ImageBuffer[24][2] ), .B(\ImageBuffer[25][2] ), .C(
        \ImageBuffer[26][2] ), .D(\ImageBuffer[27][2] ), .S0(n3346), .S1(n3485), .Y(n4530) );
  MX4X1 U5093 ( .A(\ImageBuffer[12][2] ), .B(\ImageBuffer[13][2] ), .C(
        \ImageBuffer[14][2] ), .D(\ImageBuffer[15][2] ), .S0(n3347), .S1(n3484), .Y(n4534) );
  MX4XL U5094 ( .A(\ImageBuffer[28][2] ), .B(\ImageBuffer[29][2] ), .C(
        \ImageBuffer[30][2] ), .D(\ImageBuffer[31][2] ), .S0(n3506), .S1(n3482), .Y(n4529) );
  MX4XL U5095 ( .A(\ImageBuffer[20][2] ), .B(\ImageBuffer[21][2] ), .C(
        \ImageBuffer[22][2] ), .D(\ImageBuffer[23][2] ), .S0(n3342), .S1(n3483), .Y(n4531) );
  INVX4 U5096 ( .A(n7488), .Y(n5606) );
  INVX1 U5097 ( .A(n7956), .Y(n5941) );
  INVX1 U5098 ( .A(n7959), .Y(n5940) );
  OR3X2 U5099 ( .A(n5154), .B(n5153), .C(n5152), .Y(n3569) );
  NAND3X2 U5100 ( .A(N2696), .B(N2695), .C(N2697), .Y(n8075) );
  NAND3X6 U5101 ( .A(N2707), .B(N2706), .C(N2708), .Y(n8074) );
  NOR2X1 U5102 ( .A(n5284), .B(n5296), .Y(n5297) );
  BUFX16 U5103 ( .A(n3479), .Y(n5124) );
  OAI21X1 U5104 ( .A0(n5067), .A1(n4908), .B0(n7568), .Y(n7561) );
  OAI21X1 U5105 ( .A0(n5065), .A1(n4908), .B0(n7545), .Y(n7538) );
  OAI21X1 U5106 ( .A0(n5065), .A1(n4890), .B0(n7342), .Y(n7335) );
  OAI21X1 U5107 ( .A0(n3558), .A1(n4890), .B0(n7412), .Y(n7403) );
  OAI21X1 U5108 ( .A0(n5071), .A1(n4908), .B0(n7614), .Y(n7606) );
  OAI21X1 U5109 ( .A0(n5069), .A1(n7935), .B0(n7997), .Y(n7990) );
  OAI21X1 U5110 ( .A0(n5070), .A1(n4908), .B0(n7602), .Y(n7595) );
  OAI21X1 U5111 ( .A0(n5070), .A1(n4890), .B0(n7399), .Y(n7392) );
  OAI21X1 U5112 ( .A0(n5068), .A1(n4908), .B0(n7579), .Y(n7572) );
  OAI21X1 U5113 ( .A0(n5068), .A1(n4890), .B0(n7376), .Y(n7369) );
  OAI21X1 U5114 ( .A0(n5067), .A1(n4890), .B0(n7365), .Y(n7358) );
  NOR2X1 U5115 ( .A(n5277), .B(n4865), .Y(n5235) );
  OAI2BB1XL U5116 ( .A0N(n5324), .A1N(n5077), .B0(n4866), .Y(n5323) );
  NOR2XL U5117 ( .A(n5103), .B(N2766), .Y(n5397) );
  OAI21X1 U5118 ( .A0(n5070), .A1(n4899), .B0(n7499), .Y(n7492) );
  OAI21X1 U5119 ( .A0(n5068), .A1(n4899), .B0(n7476), .Y(n7469) );
  OAI21X1 U5120 ( .A0(n5067), .A1(n4899), .B0(n7465), .Y(n7458) );
  OAI21X1 U5121 ( .A0(n5065), .A1(n4899), .B0(n7442), .Y(n7435) );
  OAI21X1 U5122 ( .A0(n4881), .A1(n5070), .B0(n7290), .Y(n7283) );
  OAI21X1 U5123 ( .A0(n4881), .A1(n5068), .B0(n7263), .Y(n7256) );
  OAI21X1 U5124 ( .A0(n4881), .A1(n5067), .B0(n7248), .Y(n7241) );
  OAI21X1 U5125 ( .A0(n4881), .A1(n5065), .B0(n7218), .Y(n7211) );
  OAI21X1 U5126 ( .A0(n5071), .A1(n4899), .B0(n7513), .Y(n7503) );
  OAI21X1 U5127 ( .A0(n4881), .A1(n5071), .B0(n7305), .Y(n7296) );
  OAI21X1 U5128 ( .A0(n4881), .A1(n5069), .B0(n7275), .Y(n7268) );
  OAI21X1 U5129 ( .A0(n4881), .A1(n5066), .B0(n7232), .Y(n7225) );
  CLKINVX2 U5130 ( .A(n8014), .Y(n5988) );
  NAND2BXL U5131 ( .AN(n3944), .B(n4872), .Y(n5262) );
  MX4XL U5132 ( .A(n4538), .B(n4528), .C(n4533), .D(n4523), .S0(N2516), .S1(
        N2515), .Y(N2755) );
  MX4X1 U5133 ( .A(n4066), .B(n4064), .C(n4065), .D(n4063), .S0(n4109), .S1(
        n4136), .Y(n4067) );
  MX4X4 U5134 ( .A(n3706), .B(n3704), .C(n3705), .D(n3703), .S0(n3734), .S1(
        n3759), .Y(n3707) );
  MX4XL U5135 ( .A(\ImageBuffer[4][0] ), .B(\ImageBuffer[5][0] ), .C(
        \ImageBuffer[6][0] ), .D(\ImageBuffer[7][0] ), .S0(n3735), .S1(n3757), 
        .Y(n3965) );
  MX4XL U5136 ( .A(\ImageBuffer[48][7] ), .B(\ImageBuffer[49][7] ), .C(
        \ImageBuffer[50][7] ), .D(\ImageBuffer[51][7] ), .S0(n4119), .S1(n4125), .Y(n4091) );
  MX4XL U5137 ( .A(\ImageBuffer[52][1] ), .B(\ImageBuffer[53][1] ), .C(
        \ImageBuffer[54][1] ), .D(\ImageBuffer[55][1] ), .S0(n3513), .S1(n3472), .Y(n4341) );
  MX4XL U5138 ( .A(\ImageBuffer[36][7] ), .B(\ImageBuffer[37][7] ), .C(
        \ImageBuffer[38][7] ), .D(\ImageBuffer[39][7] ), .S0(n4119), .S1(n5116), .Y(n4095) );
  INVX12 U5139 ( .A(cmd[0]), .Y(n5404) );
  CLKINVX2 U5140 ( .A(n8015), .Y(n5987) );
  NAND2BXL U5141 ( .AN(N2771), .B(n3944), .Y(n5383) );
  NAND2BXL U5142 ( .AN(n3944), .B(N2771), .Y(n5373) );
  NAND4X1 U5143 ( .A(N2703), .B(N2702), .C(N2701), .D(n8075), .Y(n8066) );
  CLKINVX1 U5144 ( .A(n7865), .Y(n7862) );
  CLKINVX1 U5145 ( .A(n7842), .Y(n7839) );
  INVX1 U5146 ( .A(n8005), .Y(n5977) );
  INVX3 U5147 ( .A(n7631), .Y(n5705) );
  NAND2XL U5148 ( .A(n7532), .B(n3392), .Y(n7599) );
  NAND2XL U5149 ( .A(n7532), .B(n3395), .Y(n7576) );
  NAND2XL U5150 ( .A(n7429), .B(n3392), .Y(n7496) );
  NAND2XL U5151 ( .A(n7429), .B(n3395), .Y(n7473) );
  NAND2XL U5152 ( .A(n7329), .B(n3392), .Y(n7396) );
  NAND2XL U5153 ( .A(n7329), .B(n3395), .Y(n7373) );
  NAND2XL U5154 ( .A(n7532), .B(n7234), .Y(n7553) );
  NAND2XL U5155 ( .A(n7532), .B(n7200), .Y(n7525) );
  NAND2XL U5156 ( .A(n7429), .B(n7234), .Y(n7450) );
  NAND2XL U5157 ( .A(n7429), .B(n7200), .Y(n7423) );
  NAND2XL U5158 ( .A(n7329), .B(n7234), .Y(n7350) );
  NAND2XL U5159 ( .A(n7329), .B(n7200), .Y(n7322) );
  NAND2XL U5160 ( .A(n7234), .B(n7201), .Y(n7229) );
  NAND2XL U5161 ( .A(n7200), .B(n7201), .Y(n7191) );
  NAND2XL U5162 ( .A(n3392), .B(n7201), .Y(n7287) );
  NAND2XL U5163 ( .A(n3395), .B(n7201), .Y(n7260) );
  NAND2X2 U5164 ( .A(n3569), .B(n5151), .Y(N2695) );
  NOR2X1 U5165 ( .A(n3492), .B(n5357), .Y(n5358) );
  NOR2X1 U5166 ( .A(n5250), .B(n5101), .Y(n5275) );
  AND2X2 U5167 ( .A(n5315), .B(n5325), .Y(n5322) );
  OAI21X1 U5168 ( .A0(n5068), .A1(n4926), .B0(n7780), .Y(n7773) );
  OAI21X1 U5169 ( .A0(n5071), .A1(n7935), .B0(n8027), .Y(n8016) );
  OAI21X1 U5170 ( .A0(n5066), .A1(n7935), .B0(n7960), .Y(n7952) );
  OAI21X1 U5171 ( .A0(n3548), .A1(n7935), .B0(n7932), .Y(n7920) );
  OAI21X1 U5172 ( .A0(n5070), .A1(n4926), .B0(n7803), .Y(n7796) );
  OAI21X1 U5173 ( .A0(n5067), .A1(n4926), .B0(n7769), .Y(n7762) );
  OAI21X1 U5174 ( .A0(n5065), .A1(n4926), .B0(n7746), .Y(n7739) );
  OAI21X1 U5175 ( .A0(n5071), .A1(n4926), .B0(n7815), .Y(n7807) );
  NAND2XL U5176 ( .A(n7834), .B(n3393), .Y(n7902) );
  NAND2XL U5177 ( .A(n7834), .B(n3397), .Y(n7879) );
  NAND2XL U5178 ( .A(n7834), .B(n7250), .Y(n7868) );
  NAND2XL U5179 ( .A(n7834), .B(n3396), .Y(n7845) );
  NAND2XL U5180 ( .A(n7936), .B(n3393), .Y(n8009) );
  NAND2XL U5181 ( .A(n7936), .B(n3397), .Y(n7986) );
  NAND2XL U5182 ( .A(n7936), .B(n7250), .Y(n7974) );
  NAND2XL U5183 ( .A(n7936), .B(n3396), .Y(n7948) );
  INVX3 U5184 ( .A(n7996), .Y(n5967) );
  NAND2X2 U5185 ( .A(n5043), .B(n5411), .Y(n5408) );
  NAND2X2 U5186 ( .A(n5043), .B(n4939), .Y(n5952) );
  NAND2X2 U5187 ( .A(n5043), .B(n4938), .Y(n5943) );
  NAND2X2 U5188 ( .A(n5043), .B(n4935), .Y(n5916) );
  NAND2XL U5189 ( .A(n7429), .B(n3394), .Y(n7509) );
  NAND2XL U5190 ( .A(n7329), .B(n3394), .Y(n7408) );
  NAND2XL U5191 ( .A(n7532), .B(n3394), .Y(n7610) );
  NAND2XL U5192 ( .A(n7532), .B(n7249), .Y(n7565) );
  NAND2XL U5193 ( .A(n7532), .B(n7219), .Y(n7542) );
  NAND2XL U5194 ( .A(n7429), .B(n7249), .Y(n7462) );
  NAND2XL U5195 ( .A(n7429), .B(n7219), .Y(n7439) );
  NAND2XL U5196 ( .A(n7329), .B(n7249), .Y(n7362) );
  NAND2XL U5197 ( .A(n7329), .B(n7219), .Y(n7339) );
  NAND2XL U5198 ( .A(n7532), .B(n3391), .Y(n7587) );
  NAND2XL U5199 ( .A(n7429), .B(n3391), .Y(n7484) );
  NAND2XL U5200 ( .A(n7329), .B(n3391), .Y(n7384) );
  NAND2XL U5201 ( .A(n3391), .B(n7201), .Y(n7272) );
  NAND2XL U5202 ( .A(n7249), .B(n7201), .Y(n7245) );
  NAND2XL U5203 ( .A(n7219), .B(n7201), .Y(n7215) );
  NAND2XL U5204 ( .A(n3394), .B(n7201), .Y(n7300) );
  NAND2X4 U5205 ( .A(n3523), .B(n8063), .Y(n8072) );
  CLKINVX1 U5206 ( .A(n4865), .Y(n5186) );
  INVX1 U5207 ( .A(n4865), .Y(n5156) );
  OAI2BB1XL U5208 ( .A0N(n5353), .A1N(n5077), .B0(n4873), .Y(n5352) );
  OAI21X1 U5209 ( .A0(n5071), .A1(n7833), .B0(n7914), .Y(n7906) );
  OAI21X1 U5210 ( .A0(n5070), .A1(n7833), .B0(n7902), .Y(n7895) );
  OAI21X1 U5211 ( .A0(n5068), .A1(n7833), .B0(n7879), .Y(n7872) );
  OAI21X1 U5212 ( .A0(n5065), .A1(n4917), .B0(n7645), .Y(n7638) );
  OAI21X1 U5213 ( .A0(n5070), .A1(n4917), .B0(n7702), .Y(n7695) );
  OAI21X1 U5214 ( .A0(n5068), .A1(n4917), .B0(n7679), .Y(n7672) );
  OAI21X1 U5215 ( .A0(n5067), .A1(n4917), .B0(n7668), .Y(n7661) );
  OAI21X1 U5216 ( .A0(n5067), .A1(n7833), .B0(n7868), .Y(n7861) );
  OAI21X1 U5217 ( .A0(n5065), .A1(n7833), .B0(n7845), .Y(n7838) );
  OAI21X1 U5218 ( .A0(n5069), .A1(n7833), .B0(n7890), .Y(n7883) );
  OAI21X1 U5219 ( .A0(n5066), .A1(n7833), .B0(n7856), .Y(n7849) );
  OAI21X1 U5220 ( .A0(n5052), .A1(n7833), .B0(n7830), .Y(n7822) );
  NAND2X2 U5221 ( .A(n5041), .B(n4887), .Y(n5529) );
  NAND2X2 U5222 ( .A(n5041), .B(n4900), .Y(n5628) );
  NAND2X2 U5223 ( .A(n5041), .B(n4896), .Y(n5601) );
  NAND2X2 U5224 ( .A(n7179), .B(n4893), .Y(n5574) );
  NAND2X2 U5225 ( .A(n5041), .B(n4891), .Y(n5556) );
  NAND2X2 U5226 ( .A(n5041), .B(n4894), .Y(n5583) );
  NAND2X2 U5227 ( .A(n5041), .B(n4892), .Y(n5565) );
  NAND2X2 U5228 ( .A(n5041), .B(n4897), .Y(n5610) );
  NAND2X2 U5229 ( .A(n5042), .B(n4903), .Y(n5655) );
  NAND2X2 U5230 ( .A(n5041), .B(n4895), .Y(n5592) );
  NAND2X2 U5231 ( .A(n5042), .B(n4906), .Y(n5682) );
  NAND2X2 U5232 ( .A(n5042), .B(n4904), .Y(n5664) );
  NAND2X2 U5233 ( .A(n5041), .B(n4888), .Y(n5538) );
  NAND2X2 U5234 ( .A(n5044), .B(n4886), .Y(n5520) );
  NAND2X2 U5235 ( .A(n5044), .B(n4883), .Y(n5493) );
  NAND2X2 U5236 ( .A(n5042), .B(n4907), .Y(n5691) );
  NAND2X2 U5237 ( .A(n5042), .B(n4910), .Y(n5709) );
  NAND2X2 U5238 ( .A(n5042), .B(n4913), .Y(n5736) );
  NAND2X2 U5239 ( .A(n5041), .B(n4898), .Y(n5619) );
  NAND2X2 U5240 ( .A(n5044), .B(n4889), .Y(n5547) );
  NAND2X2 U5241 ( .A(n5044), .B(n4922), .Y(n5808) );
  NAND2X2 U5242 ( .A(n5044), .B(n4921), .Y(n5799) );
  NAND2X2 U5243 ( .A(n5043), .B(n4941), .Y(n5970) );
  NAND2X2 U5244 ( .A(n5043), .B(n4937), .Y(n5934) );
  NAND2X2 U5245 ( .A(n5043), .B(n4936), .Y(n5925) );
  NAND2X2 U5246 ( .A(n5043), .B(n4934), .Y(n5907) );
  NAND2X2 U5247 ( .A(n5043), .B(n4932), .Y(n5889) );
  NAND2X2 U5248 ( .A(n5043), .B(n4940), .Y(n5961) );
  NAND2X2 U5249 ( .A(n5043), .B(n4933), .Y(n5898) );
  NAND2X2 U5250 ( .A(n5043), .B(n4931), .Y(n5880) );
  NAND3XL U5251 ( .A(n3755), .B(n3939), .C(N2495), .Y(n3547) );
  MX4X2 U5252 ( .A(n4578), .B(n4568), .C(n4573), .D(n4563), .S0(N2516), .S1(
        N2515), .Y(N2753) );
  AOI222X2 U5253 ( .A0(N2744), .A1(n4943), .B0(sum[7]), .B1(n5987), .C0(N2752), 
        .C1(n5988), .Y(n6385) );
  NAND2X2 U5254 ( .A(N2742), .B(n4943), .Y(n3563) );
  NAND2X6 U5255 ( .A(sum[9]), .B(n5987), .Y(n3564) );
  NAND2X2 U5256 ( .A(N2750), .B(n5988), .Y(n3565) );
  MX4X1 U5257 ( .A(n3848), .B(n3846), .C(n3847), .D(n3845), .S0(n3933), .S1(
        n3409), .Y(n3849) );
  AO22X1 U5258 ( .A0(N2632), .A1(n3476), .B0(N2495), .B1(n3477), .Y(n8049) );
  XNOR2XL U5259 ( .A(\sub_168_aco/carry[2] ), .B(N2495), .Y(N2632) );
  XOR2XL U5260 ( .A(n5125), .B(\add_162_S2_aco/carry[4] ), .Y(N2624) );
  AO22XL U5261 ( .A0(n8037), .A1(n5104), .B0(N2570), .B1(n8038), .Y(n3329) );
  AO22XL U5262 ( .A0(n8037), .A1(N2519), .B0(N2569), .B1(n8038), .Y(n3330) );
  AO22XL U5263 ( .A0(n8037), .A1(n5105), .B0(N2568), .B1(n8038), .Y(n3331) );
  AO22XL U5264 ( .A0(n8037), .A1(n5106), .B0(n5107), .B1(n8038), .Y(n3332) );
  OAI21XL U5265 ( .A0(n6580), .A1(n5979), .B0(n6581), .Y(n8345) );
  OAI21XL U5266 ( .A0(n6382), .A1(n5979), .B0(n6383), .Y(n8281) );
  MX4XL U5267 ( .A(\ImageBuffer[12][0] ), .B(\ImageBuffer[13][0] ), .C(
        \ImageBuffer[14][0] ), .D(\ImageBuffer[15][0] ), .S0(n3735), .S1(n5116), .Y(n3963) );
  MX4X1 U5268 ( .A(\ImageBuffer[16][0] ), .B(\ImageBuffer[17][0] ), .C(
        \ImageBuffer[18][0] ), .D(\ImageBuffer[19][0] ), .S0(n3343), .S1(n3485), .Y(n4492) );
  MX4X1 U5269 ( .A(\ImageBuffer[60][3] ), .B(\ImageBuffer[61][3] ), .C(
        \ImageBuffer[62][3] ), .D(\ImageBuffer[63][3] ), .S0(n3741), .S1(n4126), .Y(n3633) );
  MX4X1 U5270 ( .A(\ImageBuffer[56][3] ), .B(\ImageBuffer[57][3] ), .C(
        \ImageBuffer[58][3] ), .D(\ImageBuffer[59][3] ), .S0(n3741), .S1(n3747), .Y(n3634) );
  MX4X1 U5271 ( .A(\ImageBuffer[36][3] ), .B(\ImageBuffer[37][3] ), .C(
        \ImageBuffer[38][3] ), .D(\ImageBuffer[39][3] ), .S0(n4116), .S1(n3750), .Y(n4015) );
  MX4X1 U5272 ( .A(\ImageBuffer[44][2] ), .B(\ImageBuffer[45][2] ), .C(
        \ImageBuffer[46][2] ), .D(\ImageBuffer[47][2] ), .S0(n5120), .S1(n3921), .Y(n3805) );
  MX4X1 U5273 ( .A(n4175), .B(n4173), .C(n4174), .D(n4172), .S0(n5108), .S1(
        n3487), .Y(n4176) );
  MX4XL U5274 ( .A(\ImageBuffer[28][1] ), .B(\ImageBuffer[29][1] ), .C(
        \ImageBuffer[30][1] ), .D(\ImageBuffer[31][1] ), .S0(n3512), .S1(n3473), .Y(n4349) );
  MX4XL U5275 ( .A(\ImageBuffer[60][1] ), .B(\ImageBuffer[61][1] ), .C(
        \ImageBuffer[62][1] ), .D(\ImageBuffer[63][1] ), .S0(n3511), .S1(n3472), .Y(n4339) );
  MX4XL U5276 ( .A(\ImageBuffer[24][7] ), .B(\ImageBuffer[25][7] ), .C(
        \ImageBuffer[26][7] ), .D(\ImageBuffer[27][7] ), .S0(n3938), .S1(n3920), .Y(n3911) );
  MX4XL U5277 ( .A(\ImageBuffer[28][7] ), .B(\ImageBuffer[29][7] ), .C(
        \ImageBuffer[30][7] ), .D(\ImageBuffer[31][7] ), .S0(n4119), .S1(n3757), .Y(n4098) );
  MX4XL U5278 ( .A(n4051), .B(n4049), .C(n4050), .D(n4048), .S0(n4109), .S1(
        n4136), .Y(n4052) );
  AO22XL U5279 ( .A0(n8037), .A1(N2522), .B0(N2572), .B1(n8038), .Y(n3327) );
  AO22XL U5280 ( .A0(n8037), .A1(N2521), .B0(N2571), .B1(n8038), .Y(n3328) );
  XOR2XL U5281 ( .A(\add_122/carry[5] ), .B(IROM_A[5]), .Y(N2549) );
  NAND2X8 U5282 ( .A(n8086), .B(n8087), .Y(n8077) );
  INVXL U5283 ( .A(n7556), .Y(n7554) );
  INVXL U5284 ( .A(n7530), .Y(n7527) );
  INVXL U5285 ( .A(n7453), .Y(n7451) );
  INVXL U5286 ( .A(n7427), .Y(n7424) );
  INVXL U5287 ( .A(n7353), .Y(n7351) );
  INVXL U5288 ( .A(n7327), .Y(n7324) );
  INVXL U5289 ( .A(n7198), .Y(n7194) );
  NAND2BX2 U5290 ( .AN(n5274), .B(n5257), .Y(n5269) );
  INVX3 U5291 ( .A(n7816), .Y(n5840) );
  INVX3 U5292 ( .A(n7341), .Y(n5498) );
  OAI32XL U5293 ( .A0(n7335), .A1(n5054), .A2(n7336), .B0(n3352), .B1(n7342), 
        .Y(n7341) );
  OAI32XL U5294 ( .A0(n7990), .A1(n5059), .A2(n7991), .B0(n3351), .B1(n7997), 
        .Y(n7998) );
  NAND2XL U5295 ( .A(n3393), .B(n7204), .Y(n7290) );
  NAND2XL U5296 ( .A(n3397), .B(n7204), .Y(n7263) );
  INVXL U5297 ( .A(n7791), .Y(n7789) );
  INVXL U5298 ( .A(n7757), .Y(n7755) );
  INVXL U5299 ( .A(n7731), .Y(n7728) );
  INVXL U5300 ( .A(n7690), .Y(n7688) );
  INVXL U5301 ( .A(n7656), .Y(n7654) );
  INVXL U5302 ( .A(n7630), .Y(n7627) );
  INVXL U5303 ( .A(n7590), .Y(n7588) );
  INVXL U5304 ( .A(n7487), .Y(n7485) );
  INVXL U5305 ( .A(n7387), .Y(n7385) );
  BUFX20 U5306 ( .A(n3376), .Y(n5072) );
  OAI31X2 U5307 ( .A0(n5368), .A1(n5367), .A2(n5366), .B0(n5365), .Y(N2707) );
  NOR2X2 U5308 ( .A(n5316), .B(n5328), .Y(n5329) );
  NAND2BX2 U5309 ( .AN(n5306), .B(n5288), .Y(n5301) );
  NAND2BX2 U5310 ( .AN(n5367), .B(n5349), .Y(n5362) );
  NOR3BX1 U5311 ( .AN(n5149), .B(n5148), .C(n5134), .Y(n5135) );
  NAND2BX2 U5312 ( .AN(n5153), .B(n5136), .Y(n5148) );
  AND2X4 U5313 ( .A(n5344), .B(n5354), .Y(n5351) );
  INVX3 U5314 ( .A(n5229), .Y(N2673) );
  NOR3BX2 U5315 ( .AN(n5241), .B(n5240), .C(n5226), .Y(n5227) );
  INVX3 U5316 ( .A(n5258), .Y(N2674) );
  CLKINVX4 U5317 ( .A(n5197), .Y(n5220) );
  AOI31X2 U5318 ( .A0(n5220), .A1(n5198), .A2(n5214), .B0(n5217), .Y(n5199) );
  AOI31X2 U5319 ( .A0(n5311), .A1(n5288), .A2(n5304), .B0(n5307), .Y(n5289) );
  NAND2BX2 U5320 ( .AN(n5338), .B(n5320), .Y(n5333) );
  INVX3 U5321 ( .A(n7710), .Y(n5770) );
  NAND2XL U5322 ( .A(n7934), .B(n3394), .Y(n8023) );
  NAND2XL U5323 ( .A(n7733), .B(n3394), .Y(n7811) );
  NAND2XL U5324 ( .A(n7250), .B(n7204), .Y(n7248) );
  NAND2XL U5325 ( .A(n3396), .B(n7204), .Y(n7218) );
  INVX1 U5326 ( .A(N2497), .Y(n7515) );
  CLKINVX6 U5327 ( .A(n5078), .Y(n5076) );
  OAI211X1 U5328 ( .A0(n4866), .A1(n5202), .B0(n5201), .C0(n5200), .Y(n5204)
         );
  NOR2XL U5329 ( .A(n5085), .B(n4865), .Y(n5327) );
  NAND2BXL U5330 ( .AN(n4863), .B(n5093), .Y(n5334) );
  NAND2BXL U5331 ( .AN(N2768), .B(n3360), .Y(n5392) );
  NAND2XL U5332 ( .A(N2767), .B(n5098), .Y(n5378) );
  NAND2BXL U5333 ( .AN(n4863), .B(n4869), .Y(n5241) );
  NAND2BXL U5334 ( .AN(N2768), .B(n4869), .Y(n5302) );
  NAND2XL U5335 ( .A(n4865), .B(n5088), .Y(n5330) );
  CLKBUFX2 U5336 ( .A(n5088), .Y(n5087) );
  CLKBUFX2 U5337 ( .A(n5088), .Y(n5086) );
  NOR2XL U5338 ( .A(n5103), .B(n4861), .Y(n5339) );
  NAND2XL U5339 ( .A(N2766), .B(n5102), .Y(n5394) );
  CLKBUFX2 U5340 ( .A(n5103), .Y(n5102) );
  OAI21X1 U5341 ( .A0(n3558), .A1(n4917), .B0(n7715), .Y(n7706) );
  INVX1 U5342 ( .A(N2498), .Y(n7717) );
  NAND3XL U5343 ( .A(N2498), .B(N2497), .C(n5127), .Y(n7330) );
  MX4X2 U5344 ( .A(n4358), .B(n4348), .C(n4353), .D(n4343), .S0(N2510), .S1(
        N2509), .Y(N2748) );
  MX4X2 U5345 ( .A(n3808), .B(n3806), .C(n3807), .D(n3805), .S0(n3933), .S1(
        N2489), .Y(n3809) );
  MX4X2 U5346 ( .A(n3818), .B(n3816), .C(n3817), .D(n3815), .S0(n3933), .S1(
        N2489), .Y(n3819) );
  MX4XL U5347 ( .A(n4637), .B(n4635), .C(n4636), .D(n4634), .S0(n3496), .S1(
        n4640), .Y(n4638) );
  MX4XL U5348 ( .A(n4627), .B(n4625), .C(n4626), .D(n4624), .S0(n3496), .S1(
        n4640), .Y(n4628) );
  MX4XL U5349 ( .A(n4622), .B(n4620), .C(n4621), .D(n4619), .S0(n3496), .S1(
        n4640), .Y(n4623) );
  MX4XL U5350 ( .A(n4638), .B(n4628), .C(n4633), .D(n4623), .S0(N2516), .S1(
        N2515), .Y(N2750) );
  MX4XL U5351 ( .A(n4617), .B(n4615), .C(n4616), .D(n4614), .S0(n3496), .S1(
        n4640), .Y(n4618) );
  MX4XL U5352 ( .A(n4607), .B(n4605), .C(n4606), .D(n4604), .S0(n3496), .S1(
        n4640), .Y(n4608) );
  MX4XL U5353 ( .A(n4602), .B(n4600), .C(n4601), .D(n4599), .S0(n3496), .S1(
        n4640), .Y(n4603) );
  MX4XL U5354 ( .A(n4618), .B(n4608), .C(n4613), .D(n4603), .S0(N2516), .S1(
        N2515), .Y(N2751) );
  BUFX12 U5355 ( .A(N2761), .Y(n4870) );
  MXI4X4 U5356 ( .A(n4007), .B(n3997), .C(n4002), .D(n3992), .S0(N2498), .S1(
        N2497), .Y(n3550) );
  MXI4X4 U5357 ( .A(n3587), .B(n3577), .C(n3592), .D(n3582), .S0(n4946), .S1(
        n5126), .Y(n3551) );
  MXI4X4 U5358 ( .A(n3632), .B(n3622), .C(n3627), .D(n3617), .S0(n4946), .S1(
        n5125), .Y(n3552) );
  MX4XL U5359 ( .A(n3918), .B(n3916), .C(n3917), .D(n3915), .S0(n3933), .S1(
        n3409), .Y(n3919) );
  MX4XL U5360 ( .A(n3908), .B(n3906), .C(n3907), .D(n3905), .S0(N2490), .S1(
        n3409), .Y(n3909) );
  BUFX8 U5361 ( .A(N2759), .Y(n4868) );
  MX4X2 U5362 ( .A(n3899), .B(n3889), .C(n3894), .D(n3884), .S0(N2492), .S1(
        N2491), .Y(N2759) );
  MX4XL U5363 ( .A(n3898), .B(n3896), .C(n3897), .D(n3895), .S0(n3933), .S1(
        n3409), .Y(n3899) );
  MX4XL U5364 ( .A(n3888), .B(n3886), .C(n3887), .D(n3885), .S0(n3933), .S1(
        n3409), .Y(n3889) );
  MX4XL U5365 ( .A(n3863), .B(n3861), .C(n3862), .D(n3860), .S0(n3933), .S1(
        n3409), .Y(n3864) );
  MX4XL U5366 ( .A(n3868), .B(n3866), .C(n3867), .D(n3865), .S0(n3933), .S1(
        n3409), .Y(n3869) );
  MX4X4 U5367 ( .A(n3712), .B(n3702), .C(n3707), .D(n3697), .S0(n4946), .S1(
        n5125), .Y(N2775) );
  MX4XL U5368 ( .A(n3696), .B(n3694), .C(n3695), .D(n3693), .S0(n3734), .S1(
        n3759), .Y(n3697) );
  MX4X2 U5369 ( .A(n4558), .B(n4548), .C(n4553), .D(n4543), .S0(N2516), .S1(
        N2515), .Y(N2754) );
  MX4XL U5370 ( .A(n4467), .B(n4465), .C(n4466), .D(n4464), .S0(n3503), .S1(
        n3495), .Y(n4468) );
  MX4XL U5371 ( .A(n4462), .B(n4460), .C(n4461), .D(n4459), .S0(n3503), .S1(
        n3495), .Y(n4463) );
  MX4XL U5372 ( .A(n4458), .B(n4448), .C(n4453), .D(n4443), .S0(N2510), .S1(
        N2509), .Y(N2743) );
  MX4XL U5373 ( .A(n4457), .B(n4455), .C(n4456), .D(n4454), .S0(n3503), .S1(
        n3495), .Y(n4458) );
  MX4XL U5374 ( .A(n4447), .B(n4445), .C(n4446), .D(n4444), .S0(n3503), .S1(
        n3495), .Y(n4448) );
  MX4XL U5375 ( .A(n4442), .B(n4440), .C(n4441), .D(n4439), .S0(n3503), .S1(
        n3495), .Y(n4443) );
  MXI4X4 U5376 ( .A(n3953), .B(n3951), .C(n3952), .D(n3950), .S0(n4109), .S1(
        n3758), .Y(n3556) );
  MX4XL U5377 ( .A(n4280), .B(n4278), .C(n4279), .D(n4277), .S0(n5108), .S1(
        n3487), .Y(n4281) );
  MX4XL U5378 ( .A(n4285), .B(n4283), .C(n4284), .D(n4282), .S0(n5108), .S1(
        n3487), .Y(n4286) );
  MX4XL U5379 ( .A(n4295), .B(n4293), .C(n4294), .D(n4292), .S0(n5108), .S1(
        n3487), .Y(n4296) );
  MX4XL U5380 ( .A(n4245), .B(n4243), .C(n4244), .D(n4242), .S0(n5108), .S1(
        n3487), .Y(n4246) );
  MX4XL U5381 ( .A(n4240), .B(n4238), .C(n4239), .D(n4237), .S0(n5108), .S1(
        n3487), .Y(n4241) );
  MX4XL U5382 ( .A(n4250), .B(n4248), .C(n4249), .D(n4247), .S0(n5108), .S1(
        n3487), .Y(n4251) );
  BUFX8 U5383 ( .A(N2774), .Y(n4861) );
  MX4XL U5384 ( .A(n3731), .B(n3729), .C(n3730), .D(n3728), .S0(n3734), .S1(
        n3759), .Y(n3732) );
  MX4XL U5385 ( .A(n3721), .B(n3719), .C(n3720), .D(n3718), .S0(n3734), .S1(
        n3759), .Y(n3722) );
  MX4XL U5386 ( .A(n4056), .B(n4054), .C(n4055), .D(n4053), .S0(n4109), .S1(
        n4136), .Y(n4057) );
  AO22XL U5387 ( .A0(N2634), .A1(n3476), .B0(N2614), .B1(n3477), .Y(n8053) );
  NAND3XL U5388 ( .A(N2497), .B(n5128), .C(N2498), .Y(n7202) );
  NAND2X1 U5389 ( .A(n7922), .B(n5115), .Y(n3560) );
  CLKBUFX2 U5390 ( .A(n5121), .Y(n5120) );
  NOR2XL U5391 ( .A(n5400), .B(n8061), .Y(N2541) );
  OR2XL U5392 ( .A(n5125), .B(\sub_168_aco/carry[4] ), .Y(
        \sub_168_aco/carry[5] ) );
  OR2XL U5393 ( .A(n5125), .B(\sub_157_S2_aco/carry[4] ), .Y(
        \sub_157_S2_aco/carry[5] ) );
  CLKINVX1 U5394 ( .A(n5107), .Y(n5106) );
  MXI2XL U5395 ( .A(\ImageBuffer[30][4] ), .B(n4988), .S0(n4910), .Y(n6491) );
  MXI2XL U5396 ( .A(\ImageBuffer[33][4] ), .B(n4987), .S0(n4906), .Y(n6482) );
  MXI2XL U5397 ( .A(\ImageBuffer[35][4] ), .B(n4988), .S0(n4904), .Y(n6476) );
  MXI2XL U5398 ( .A(\ImageBuffer[36][4] ), .B(n4988), .S0(n4903), .Y(n6473) );
  MXI2XL U5399 ( .A(\ImageBuffer[38][4] ), .B(n4988), .S0(n4901), .Y(n6467) );
  MXI2XL U5400 ( .A(\ImageBuffer[41][4] ), .B(n4988), .S0(n4897), .Y(n6458) );
  MXI2XL U5401 ( .A(\ImageBuffer[43][4] ), .B(n4988), .S0(n4895), .Y(n6452) );
  MXI2XL U5402 ( .A(\ImageBuffer[14][4] ), .B(n4987), .S0(n4928), .Y(n6539) );
  MXI2XL U5403 ( .A(\ImageBuffer[13][4] ), .B(n4987), .S0(n4929), .Y(n6542) );
  MXI2XL U5404 ( .A(\ImageBuffer[15][4] ), .B(n4987), .S0(n4927), .Y(n6536) );
  MXI2XL U5405 ( .A(\ImageBuffer[18][4] ), .B(n4987), .S0(n4923), .Y(n6527) );
  MXI2XL U5406 ( .A(\ImageBuffer[21][4] ), .B(n4987), .S0(n4920), .Y(n6518) );
  MXI2XL U5407 ( .A(\ImageBuffer[23][4] ), .B(n4987), .S0(n4918), .Y(n6512) );
  MXI2XL U5408 ( .A(\ImageBuffer[26][4] ), .B(n4987), .S0(n4914), .Y(n6503) );
  MXI2XL U5409 ( .A(\ImageBuffer[29][4] ), .B(n4987), .S0(n4911), .Y(n6494) );
  MXI2XL U5410 ( .A(\ImageBuffer[31][4] ), .B(n6388), .S0(n4909), .Y(n6488) );
  MXI2XL U5411 ( .A(\ImageBuffer[34][4] ), .B(n4988), .S0(n4905), .Y(n6479) );
  MXI2XL U5412 ( .A(\ImageBuffer[37][4] ), .B(n4988), .S0(n4902), .Y(n6470) );
  MXI2XL U5413 ( .A(\ImageBuffer[39][4] ), .B(n4988), .S0(n4900), .Y(n6464) );
  MXI2XL U5414 ( .A(\ImageBuffer[42][4] ), .B(n4988), .S0(n4896), .Y(n6455) );
  MXI2XL U5415 ( .A(\ImageBuffer[45][4] ), .B(n4988), .S0(n4893), .Y(n6446) );
  MXI2XL U5416 ( .A(\ImageBuffer[47][4] ), .B(n4988), .S0(n4891), .Y(n6440) );
  MXI2XL U5417 ( .A(\ImageBuffer[50][4] ), .B(n6388), .S0(n4887), .Y(n6431) );
  MXI2XL U5418 ( .A(\ImageBuffer[53][4] ), .B(n4986), .S0(n4884), .Y(n6422) );
  MXI2XL U5419 ( .A(\ImageBuffer[55][4] ), .B(n4987), .S0(n4882), .Y(n6416) );
  MXI2XL U5420 ( .A(\ImageBuffer[56][4] ), .B(n4988), .S0(n4880), .Y(n6413) );
  MXI2XL U5421 ( .A(\ImageBuffer[17][4] ), .B(n4987), .S0(n4924), .Y(n6530) );
  MXI2XL U5422 ( .A(\ImageBuffer[20][4] ), .B(n4987), .S0(n4921), .Y(n6521) );
  MXI2XL U5423 ( .A(\ImageBuffer[22][4] ), .B(n4987), .S0(n4919), .Y(n6515) );
  MXI2XL U5424 ( .A(\ImageBuffer[24][4] ), .B(n4987), .S0(n4916), .Y(n6509) );
  MXI2XL U5425 ( .A(\ImageBuffer[40][4] ), .B(n4988), .S0(n4898), .Y(n6461) );
  MXI2XL U5426 ( .A(\ImageBuffer[48][4] ), .B(n4986), .S0(n4889), .Y(n6437) );
  MXI2XL U5427 ( .A(\ImageBuffer[57][4] ), .B(n4987), .S0(n4879), .Y(n6410) );
  MXI2XL U5428 ( .A(\ImageBuffer[59][4] ), .B(n4988), .S0(n4877), .Y(n6404) );
  MXI2XL U5429 ( .A(\ImageBuffer[25][4] ), .B(n4987), .S0(n4915), .Y(n6506) );
  MXI2XL U5430 ( .A(\ImageBuffer[27][4] ), .B(n6388), .S0(n4913), .Y(n6500) );
  MXI2XL U5431 ( .A(\ImageBuffer[28][4] ), .B(n4988), .S0(n4912), .Y(n6497) );
  MXI2XL U5432 ( .A(\ImageBuffer[49][4] ), .B(n4987), .S0(n4888), .Y(n6434) );
  MXI2XL U5433 ( .A(\ImageBuffer[51][4] ), .B(n4988), .S0(n4886), .Y(n6428) );
  MXI2XL U5434 ( .A(\ImageBuffer[52][4] ), .B(n4986), .S0(n4885), .Y(n6425) );
  MXI2XL U5435 ( .A(\ImageBuffer[54][4] ), .B(n4986), .S0(n4883), .Y(n6419) );
  MXI2XL U5436 ( .A(\ImageBuffer[32][4] ), .B(n4988), .S0(n4907), .Y(n6485) );
  MXI2XL U5437 ( .A(\ImageBuffer[12][4] ), .B(n4987), .S0(n4930), .Y(n6545) );
  MXI2XL U5438 ( .A(\ImageBuffer[9][1] ), .B(n6980), .S0(n4933), .Y(n7146) );
  MXI2XL U5439 ( .A(\ImageBuffer[11][1] ), .B(n5026), .S0(n4931), .Y(n7140) );
  MXI2XL U5440 ( .A(\ImageBuffer[30][1] ), .B(n5027), .S0(n4910), .Y(n7083) );
  MXI2XL U5441 ( .A(\ImageBuffer[33][1] ), .B(n5026), .S0(n4906), .Y(n7074) );
  MXI2XL U5442 ( .A(\ImageBuffer[35][1] ), .B(n5027), .S0(n4904), .Y(n7068) );
  MXI2XL U5443 ( .A(\ImageBuffer[36][1] ), .B(n5026), .S0(n4903), .Y(n7065) );
  MXI2XL U5444 ( .A(\ImageBuffer[38][1] ), .B(n5026), .S0(n4901), .Y(n7059) );
  MXI2XL U5445 ( .A(\ImageBuffer[41][1] ), .B(n5026), .S0(n4897), .Y(n7050) );
  MXI2XL U5446 ( .A(\ImageBuffer[43][1] ), .B(n5026), .S0(n4895), .Y(n7044) );
  MXI2XL U5447 ( .A(\ImageBuffer[2][1] ), .B(n5027), .S0(n4940), .Y(n7167) );
  MXI2XL U5448 ( .A(\ImageBuffer[14][1] ), .B(n5025), .S0(n4928), .Y(n7131) );
  MXI2XL U5449 ( .A(\ImageBuffer[5][1] ), .B(n5025), .S0(n4937), .Y(n7158) );
  MXI2XL U5450 ( .A(\ImageBuffer[7][1] ), .B(n6980), .S0(n4935), .Y(n7152) );
  MXI2XL U5451 ( .A(\ImageBuffer[10][1] ), .B(n5026), .S0(n4932), .Y(n7143) );
  MXI2XL U5452 ( .A(\ImageBuffer[13][1] ), .B(n5025), .S0(n4929), .Y(n7134) );
  MXI2XL U5453 ( .A(\ImageBuffer[15][1] ), .B(n5025), .S0(n4927), .Y(n7128) );
  MXI2XL U5454 ( .A(\ImageBuffer[18][1] ), .B(n5025), .S0(n4923), .Y(n7119) );
  MXI2XL U5455 ( .A(\ImageBuffer[21][1] ), .B(n5025), .S0(n4920), .Y(n7110) );
  MXI2XL U5456 ( .A(\ImageBuffer[23][1] ), .B(n5025), .S0(n4918), .Y(n7104) );
  MXI2XL U5457 ( .A(\ImageBuffer[26][1] ), .B(n5026), .S0(n4914), .Y(n7095) );
  MXI2XL U5458 ( .A(\ImageBuffer[29][1] ), .B(n5026), .S0(n4911), .Y(n7086) );
  MXI2XL U5459 ( .A(\ImageBuffer[31][1] ), .B(n5025), .S0(n4909), .Y(n7080) );
  MXI2XL U5460 ( .A(\ImageBuffer[34][1] ), .B(n5027), .S0(n4905), .Y(n7071) );
  MXI2XL U5461 ( .A(\ImageBuffer[37][1] ), .B(n5026), .S0(n4902), .Y(n7062) );
  MXI2XL U5462 ( .A(\ImageBuffer[39][1] ), .B(n5026), .S0(n4900), .Y(n7056) );
  MXI2XL U5463 ( .A(\ImageBuffer[42][1] ), .B(n5026), .S0(n4896), .Y(n7047) );
  MXI2XL U5464 ( .A(\ImageBuffer[45][1] ), .B(n5026), .S0(n4893), .Y(n7038) );
  MXI2XL U5465 ( .A(\ImageBuffer[47][1] ), .B(n5026), .S0(n4891), .Y(n7032) );
  MXI2XL U5466 ( .A(\ImageBuffer[53][1] ), .B(n5027), .S0(n4884), .Y(n7014) );
  MXI2XL U5467 ( .A(\ImageBuffer[55][1] ), .B(n5027), .S0(n4882), .Y(n7008) );
  MXI2XL U5468 ( .A(\ImageBuffer[1][1] ), .B(n5027), .S0(n4941), .Y(n7170) );
  MXI2XL U5469 ( .A(\ImageBuffer[3][1] ), .B(n5026), .S0(n4939), .Y(n7164) );
  MXI2XL U5470 ( .A(\ImageBuffer[4][1] ), .B(n5027), .S0(n4938), .Y(n7161) );
  MXI2XL U5471 ( .A(\ImageBuffer[6][1] ), .B(n5025), .S0(n4936), .Y(n7155) );
  MXI2XL U5472 ( .A(\ImageBuffer[17][1] ), .B(n5025), .S0(n4924), .Y(n7122) );
  MXI2XL U5473 ( .A(\ImageBuffer[20][1] ), .B(n5025), .S0(n4921), .Y(n7113) );
  MXI2XL U5474 ( .A(\ImageBuffer[22][1] ), .B(n5025), .S0(n4919), .Y(n7107) );
  MXI2XL U5475 ( .A(\ImageBuffer[24][1] ), .B(n5026), .S0(n4916), .Y(n7101) );
  MXI2XL U5476 ( .A(\ImageBuffer[40][1] ), .B(n5026), .S0(n4898), .Y(n7053) );
  MXI2XL U5477 ( .A(\ImageBuffer[48][1] ), .B(n5027), .S0(n4889), .Y(n7029) );
  MXI2XL U5478 ( .A(\ImageBuffer[57][1] ), .B(n5027), .S0(n4879), .Y(n7002) );
  MXI2XL U5479 ( .A(\ImageBuffer[59][1] ), .B(n5027), .S0(n4877), .Y(n6996) );
  MXI2XL U5480 ( .A(\ImageBuffer[25][1] ), .B(n5026), .S0(n4915), .Y(n7098) );
  MXI2XL U5481 ( .A(\ImageBuffer[27][1] ), .B(n6980), .S0(n4913), .Y(n7092) );
  MXI2XL U5482 ( .A(\ImageBuffer[28][1] ), .B(n5027), .S0(n4912), .Y(n7089) );
  MXI2XL U5483 ( .A(\ImageBuffer[49][1] ), .B(n5027), .S0(n4888), .Y(n7026) );
  MXI2XL U5484 ( .A(\ImageBuffer[51][1] ), .B(n5027), .S0(n4886), .Y(n7020) );
  MXI2XL U5485 ( .A(\ImageBuffer[52][1] ), .B(n5027), .S0(n4885), .Y(n7017) );
  MXI2XL U5486 ( .A(\ImageBuffer[54][1] ), .B(n5027), .S0(n4883), .Y(n7011) );
  MXI2XL U5487 ( .A(\ImageBuffer[32][1] ), .B(n5027), .S0(n4907), .Y(n7077) );
  MXI2XL U5488 ( .A(\ImageBuffer[12][1] ), .B(n5025), .S0(n4930), .Y(n7137) );
  MXI2XL U5489 ( .A(\ImageBuffer[19][7] ), .B(n4948), .S0(n4922), .Y(n5809) );
  MXI2XL U5490 ( .A(\ImageBuffer[30][5] ), .B(n4974), .S0(n4910), .Y(n6293) );
  MXI2XL U5491 ( .A(\ImageBuffer[30][6] ), .B(n4960), .S0(n4910), .Y(n6095) );
  MXI2XL U5492 ( .A(\ImageBuffer[30][7] ), .B(n4949), .S0(n4910), .Y(n5710) );
  MXI2XL U5493 ( .A(\ImageBuffer[33][5] ), .B(n4974), .S0(n4906), .Y(n6284) );
  MXI2XL U5494 ( .A(\ImageBuffer[33][6] ), .B(n4960), .S0(n4906), .Y(n6086) );
  MXI2XL U5495 ( .A(\ImageBuffer[33][7] ), .B(n4949), .S0(n4906), .Y(n5683) );
  MXI2XL U5496 ( .A(\ImageBuffer[35][5] ), .B(n4974), .S0(n4904), .Y(n6278) );
  MXI2XL U5497 ( .A(\ImageBuffer[35][6] ), .B(n4960), .S0(n4904), .Y(n6080) );
  MXI2XL U5498 ( .A(\ImageBuffer[35][7] ), .B(n4949), .S0(n4904), .Y(n5665) );
  MXI2XL U5499 ( .A(\ImageBuffer[36][5] ), .B(n4975), .S0(n4903), .Y(n6275) );
  MXI2XL U5500 ( .A(\ImageBuffer[38][5] ), .B(n4975), .S0(n4901), .Y(n6269) );
  MXI2XL U5501 ( .A(\ImageBuffer[38][6] ), .B(n4961), .S0(n4901), .Y(n6071) );
  MXI2XL U5502 ( .A(\ImageBuffer[43][5] ), .B(n4975), .S0(n4895), .Y(n6254) );
  MXI2XL U5503 ( .A(\ImageBuffer[43][6] ), .B(n4961), .S0(n4895), .Y(n6056) );
  MXI2XL U5504 ( .A(\ImageBuffer[14][5] ), .B(n4974), .S0(n4928), .Y(n6341) );
  MXI2XL U5505 ( .A(\ImageBuffer[14][6] ), .B(n4960), .S0(n4928), .Y(n6143) );
  MXI2XL U5506 ( .A(\ImageBuffer[14][7] ), .B(n4948), .S0(n4928), .Y(n5854) );
  MXI2XL U5507 ( .A(\ImageBuffer[13][5] ), .B(n4976), .S0(n4929), .Y(n6344) );
  MXI2XL U5508 ( .A(\ImageBuffer[13][6] ), .B(n4962), .S0(n4929), .Y(n6146) );
  MXI2XL U5509 ( .A(\ImageBuffer[13][7] ), .B(n4948), .S0(n4929), .Y(n5863) );
  MXI2XL U5510 ( .A(\ImageBuffer[15][5] ), .B(n4976), .S0(n4927), .Y(n6338) );
  MXI2XL U5511 ( .A(\ImageBuffer[15][6] ), .B(n4962), .S0(n4927), .Y(n6140) );
  MXI2XL U5512 ( .A(\ImageBuffer[15][7] ), .B(n4948), .S0(n4927), .Y(n5845) );
  MXI2XL U5513 ( .A(\ImageBuffer[18][5] ), .B(n4975), .S0(n4923), .Y(n6329) );
  MXI2XL U5514 ( .A(\ImageBuffer[18][6] ), .B(n4961), .S0(n4923), .Y(n6131) );
  MXI2XL U5515 ( .A(\ImageBuffer[18][7] ), .B(n4948), .S0(n4923), .Y(n5818) );
  MXI2XL U5516 ( .A(\ImageBuffer[21][5] ), .B(n4974), .S0(n4920), .Y(n6320) );
  MXI2XL U5517 ( .A(\ImageBuffer[21][6] ), .B(n4960), .S0(n4920), .Y(n6122) );
  MXI2XL U5518 ( .A(\ImageBuffer[21][7] ), .B(n4948), .S0(n4920), .Y(n5791) );
  MXI2XL U5519 ( .A(\ImageBuffer[23][5] ), .B(n4975), .S0(n4918), .Y(n6314) );
  MXI2XL U5520 ( .A(\ImageBuffer[23][6] ), .B(n4961), .S0(n4918), .Y(n6116) );
  MXI2XL U5521 ( .A(\ImageBuffer[23][7] ), .B(n4948), .S0(n4918), .Y(n5773) );
  MXI2XL U5522 ( .A(\ImageBuffer[26][5] ), .B(n4974), .S0(n4914), .Y(n6305) );
  MXI2XL U5523 ( .A(\ImageBuffer[26][6] ), .B(n4960), .S0(n4914), .Y(n6107) );
  MXI2XL U5524 ( .A(\ImageBuffer[26][7] ), .B(n4949), .S0(n4914), .Y(n5746) );
  MXI2XL U5525 ( .A(\ImageBuffer[29][5] ), .B(n4974), .S0(n4911), .Y(n6296) );
  MXI2XL U5526 ( .A(\ImageBuffer[29][6] ), .B(n4960), .S0(n4911), .Y(n6098) );
  MXI2XL U5527 ( .A(\ImageBuffer[29][7] ), .B(n4949), .S0(n4911), .Y(n5719) );
  MXI2XL U5528 ( .A(\ImageBuffer[31][5] ), .B(n4974), .S0(n4909), .Y(n6290) );
  MXI2XL U5529 ( .A(\ImageBuffer[31][6] ), .B(n4960), .S0(n4909), .Y(n6092) );
  MXI2XL U5530 ( .A(\ImageBuffer[31][7] ), .B(n4949), .S0(n4909), .Y(n5701) );
  MXI2XL U5531 ( .A(\ImageBuffer[34][5] ), .B(n4974), .S0(n4905), .Y(n6281) );
  MXI2XL U5532 ( .A(\ImageBuffer[34][6] ), .B(n4960), .S0(n4905), .Y(n6083) );
  MXI2XL U5533 ( .A(\ImageBuffer[34][7] ), .B(n4949), .S0(n4905), .Y(n5674) );
  MXI2XL U5534 ( .A(\ImageBuffer[37][5] ), .B(n4975), .S0(n4902), .Y(n6272) );
  MXI2XL U5535 ( .A(\ImageBuffer[37][6] ), .B(n4961), .S0(n4902), .Y(n6074) );
  MXI2XL U5536 ( .A(\ImageBuffer[37][7] ), .B(n4950), .S0(n4902), .Y(n5647) );
  MXI2XL U5537 ( .A(\ImageBuffer[39][5] ), .B(n4975), .S0(n4900), .Y(n6266) );
  MXI2XL U5538 ( .A(\ImageBuffer[39][6] ), .B(n4961), .S0(n4900), .Y(n6068) );
  MXI2XL U5539 ( .A(\ImageBuffer[39][7] ), .B(n4950), .S0(n4900), .Y(n5629) );
  MXI2XL U5540 ( .A(\ImageBuffer[42][5] ), .B(n4975), .S0(n4896), .Y(n6257) );
  MXI2XL U5541 ( .A(\ImageBuffer[42][6] ), .B(n4961), .S0(n4896), .Y(n6059) );
  MXI2XL U5542 ( .A(\ImageBuffer[42][7] ), .B(n4950), .S0(n4896), .Y(n5602) );
  MXI2XL U5543 ( .A(\ImageBuffer[45][5] ), .B(n4975), .S0(n4893), .Y(n6248) );
  MXI2XL U5544 ( .A(\ImageBuffer[45][6] ), .B(n4961), .S0(n4893), .Y(n6050) );
  MXI2XL U5545 ( .A(\ImageBuffer[45][7] ), .B(n4950), .S0(n4893), .Y(n5575) );
  MXI2XL U5546 ( .A(\ImageBuffer[47][5] ), .B(n4975), .S0(n4891), .Y(n6242) );
  MXI2XL U5547 ( .A(\ImageBuffer[47][6] ), .B(n4961), .S0(n4891), .Y(n6044) );
  MXI2XL U5548 ( .A(\ImageBuffer[47][7] ), .B(n4950), .S0(n4891), .Y(n5557) );
  MXI2XL U5549 ( .A(\ImageBuffer[50][7] ), .B(n4948), .S0(n4887), .Y(n5530) );
  MXI2XL U5550 ( .A(\ImageBuffer[53][5] ), .B(n4976), .S0(n4884), .Y(n6224) );
  MXI2XL U5551 ( .A(\ImageBuffer[53][7] ), .B(n4949), .S0(n4884), .Y(n5503) );
  MXI2XL U5552 ( .A(\ImageBuffer[55][5] ), .B(n4976), .S0(n4882), .Y(n6218) );
  MXI2XL U5553 ( .A(\ImageBuffer[55][6] ), .B(n4962), .S0(n4882), .Y(n6020) );
  MXI2XL U5554 ( .A(\ImageBuffer[55][7] ), .B(n4948), .S0(n4882), .Y(n5485) );
  MXI2XL U5555 ( .A(\ImageBuffer[56][7] ), .B(n4950), .S0(n4880), .Y(n5476) );
  MXI2XL U5556 ( .A(\ImageBuffer[58][7] ), .B(n4948), .S0(n4878), .Y(n5458) );
  MXI2XL U5557 ( .A(\ImageBuffer[17][5] ), .B(n4976), .S0(n4924), .Y(n6332) );
  MXI2XL U5558 ( .A(\ImageBuffer[17][6] ), .B(n4962), .S0(n4924), .Y(n6134) );
  MXI2XL U5559 ( .A(\ImageBuffer[17][7] ), .B(n4948), .S0(n4924), .Y(n5827) );
  MXI2XL U5560 ( .A(\ImageBuffer[20][5] ), .B(n4976), .S0(n4921), .Y(n6323) );
  MXI2XL U5561 ( .A(\ImageBuffer[20][6] ), .B(n4962), .S0(n4921), .Y(n6125) );
  MXI2XL U5562 ( .A(\ImageBuffer[20][7] ), .B(n4948), .S0(n4921), .Y(n5800) );
  MXI2XL U5563 ( .A(\ImageBuffer[22][5] ), .B(n4975), .S0(n4919), .Y(n6317) );
  MXI2XL U5564 ( .A(\ImageBuffer[22][6] ), .B(n4961), .S0(n4919), .Y(n6119) );
  MXI2XL U5565 ( .A(\ImageBuffer[22][7] ), .B(n4948), .S0(n4919), .Y(n5782) );
  MXI2XL U5566 ( .A(\ImageBuffer[24][5] ), .B(n4974), .S0(n4916), .Y(n6311) );
  MXI2XL U5567 ( .A(\ImageBuffer[24][6] ), .B(n4960), .S0(n4916), .Y(n6113) );
  MXI2XL U5568 ( .A(\ImageBuffer[24][7] ), .B(n4949), .S0(n4916), .Y(n5764) );
  MXI2XL U5569 ( .A(\ImageBuffer[40][5] ), .B(n4975), .S0(n4898), .Y(n6263) );
  MXI2XL U5570 ( .A(\ImageBuffer[40][6] ), .B(n4961), .S0(n4898), .Y(n6065) );
  MXI2XL U5571 ( .A(\ImageBuffer[40][7] ), .B(n4950), .S0(n4898), .Y(n5620) );
  MXI2XL U5572 ( .A(\ImageBuffer[48][5] ), .B(n4976), .S0(n4889), .Y(n6239) );
  MXI2XL U5573 ( .A(\ImageBuffer[48][6] ), .B(n4962), .S0(n4889), .Y(n6041) );
  MXI2XL U5574 ( .A(\ImageBuffer[48][7] ), .B(n4950), .S0(n4889), .Y(n5548) );
  MXI2XL U5575 ( .A(\ImageBuffer[57][5] ), .B(n4976), .S0(n4879), .Y(n6212) );
  MXI2XL U5576 ( .A(\ImageBuffer[57][6] ), .B(n4962), .S0(n4879), .Y(n6014) );
  MXI2XL U5577 ( .A(\ImageBuffer[57][7] ), .B(n4950), .S0(n4879), .Y(n5467) );
  MXI2XL U5578 ( .A(\ImageBuffer[59][5] ), .B(n4976), .S0(n4877), .Y(n6206) );
  MXI2XL U5579 ( .A(\ImageBuffer[59][6] ), .B(n4962), .S0(n4877), .Y(n6008) );
  MXI2XL U5580 ( .A(\ImageBuffer[59][7] ), .B(n4949), .S0(n4877), .Y(n5449) );
  MXI2XL U5581 ( .A(\ImageBuffer[25][5] ), .B(n4974), .S0(n4915), .Y(n6308) );
  MXI2XL U5582 ( .A(\ImageBuffer[25][6] ), .B(n4960), .S0(n4915), .Y(n6110) );
  MXI2XL U5583 ( .A(\ImageBuffer[25][7] ), .B(n4949), .S0(n4915), .Y(n5755) );
  MXI2XL U5584 ( .A(\ImageBuffer[27][5] ), .B(n4974), .S0(n4913), .Y(n6302) );
  MXI2XL U5585 ( .A(\ImageBuffer[27][6] ), .B(n4960), .S0(n4913), .Y(n6104) );
  MXI2XL U5586 ( .A(\ImageBuffer[27][7] ), .B(n4949), .S0(n4913), .Y(n5737) );
  MXI2XL U5587 ( .A(\ImageBuffer[28][5] ), .B(n4974), .S0(n4912), .Y(n6299) );
  MXI2XL U5588 ( .A(\ImageBuffer[28][6] ), .B(n4960), .S0(n4912), .Y(n6101) );
  MXI2XL U5589 ( .A(\ImageBuffer[28][7] ), .B(n4949), .S0(n4912), .Y(n5728) );
  MXI2XL U5590 ( .A(\ImageBuffer[49][5] ), .B(n4976), .S0(n4888), .Y(n6236) );
  MXI2XL U5591 ( .A(\ImageBuffer[49][6] ), .B(n4962), .S0(n4888), .Y(n6038) );
  MXI2XL U5592 ( .A(\ImageBuffer[49][7] ), .B(n4948), .S0(n4888), .Y(n5539) );
  MXI2XL U5593 ( .A(\ImageBuffer[51][5] ), .B(n4976), .S0(n4886), .Y(n6230) );
  MXI2XL U5594 ( .A(\ImageBuffer[51][6] ), .B(n4962), .S0(n4886), .Y(n6032) );
  MXI2XL U5595 ( .A(\ImageBuffer[51][7] ), .B(n4950), .S0(n4886), .Y(n5521) );
  MXI2XL U5596 ( .A(\ImageBuffer[52][5] ), .B(n4976), .S0(n4885), .Y(n6227) );
  MXI2XL U5597 ( .A(\ImageBuffer[52][6] ), .B(n4962), .S0(n4885), .Y(n6029) );
  MXI2XL U5598 ( .A(\ImageBuffer[52][7] ), .B(n4948), .S0(n4885), .Y(n5512) );
  MXI2XL U5599 ( .A(\ImageBuffer[54][5] ), .B(n4976), .S0(n4883), .Y(n6221) );
  MXI2XL U5600 ( .A(\ImageBuffer[54][6] ), .B(n4962), .S0(n4883), .Y(n6023) );
  MXI2XL U5601 ( .A(\ImageBuffer[54][7] ), .B(n4949), .S0(n4883), .Y(n5494) );
  MXI2XL U5602 ( .A(\ImageBuffer[32][5] ), .B(n4974), .S0(n4907), .Y(n6287) );
  MXI2XL U5603 ( .A(\ImageBuffer[32][6] ), .B(n4960), .S0(n4907), .Y(n6089) );
  MXI2XL U5604 ( .A(\ImageBuffer[32][7] ), .B(n4949), .S0(n4907), .Y(n5692) );
  MXI2XL U5605 ( .A(\ImageBuffer[12][5] ), .B(n4975), .S0(n4930), .Y(n6347) );
  MXI2XL U5606 ( .A(\ImageBuffer[12][6] ), .B(n4961), .S0(n4930), .Y(n6149) );
  MXI2XL U5607 ( .A(\ImageBuffer[12][7] ), .B(n4948), .S0(n4930), .Y(n5872) );
  MX4XL U5608 ( .A(\ImageBuffer[0][1] ), .B(\ImageBuffer[1][1] ), .C(
        \ImageBuffer[2][1] ), .D(\ImageBuffer[3][1] ), .S0(n5120), .S1(n3925), 
        .Y(n3798) );
  MX4XL U5609 ( .A(\ImageBuffer[32][1] ), .B(\ImageBuffer[33][1] ), .C(
        \ImageBuffer[34][1] ), .D(\ImageBuffer[35][1] ), .S0(n3939), .S1(n3922), .Y(n3788) );
  MX4XL U5610 ( .A(\ImageBuffer[16][7] ), .B(\ImageBuffer[17][7] ), .C(
        \ImageBuffer[18][7] ), .D(\ImageBuffer[19][7] ), .S0(n3346), .S1(n3483), .Y(n4632) );
  MX4XL U5611 ( .A(\ImageBuffer[24][7] ), .B(\ImageBuffer[25][7] ), .C(
        \ImageBuffer[26][7] ), .D(\ImageBuffer[27][7] ), .S0(n3506), .S1(n3484), .Y(n4630) );
  MX4XL U5612 ( .A(\ImageBuffer[28][7] ), .B(\ImageBuffer[29][7] ), .C(
        \ImageBuffer[30][7] ), .D(\ImageBuffer[31][7] ), .S0(n3342), .S1(n3482), .Y(n4629) );
  MX4XL U5613 ( .A(\ImageBuffer[16][6] ), .B(\ImageBuffer[17][6] ), .C(
        \ImageBuffer[18][6] ), .D(\ImageBuffer[19][6] ), .S0(n3343), .S1(n3485), .Y(n4612) );
  MX4XL U5614 ( .A(\ImageBuffer[24][6] ), .B(\ImageBuffer[25][6] ), .C(
        \ImageBuffer[26][6] ), .D(\ImageBuffer[27][6] ), .S0(n3506), .S1(n3482), .Y(n4610) );
  MX4XL U5615 ( .A(\ImageBuffer[28][6] ), .B(\ImageBuffer[29][6] ), .C(
        \ImageBuffer[30][6] ), .D(\ImageBuffer[31][6] ), .S0(n3343), .S1(n3483), .Y(n4609) );
  MX4XL U5616 ( .A(\ImageBuffer[20][1] ), .B(\ImageBuffer[21][1] ), .C(
        \ImageBuffer[22][1] ), .D(\ImageBuffer[23][1] ), .S0(n3486), .S1(n3339), .Y(n3792) );
  MX4XL U5617 ( .A(\ImageBuffer[4][1] ), .B(\ImageBuffer[5][1] ), .C(
        \ImageBuffer[6][1] ), .D(\ImageBuffer[7][1] ), .S0(n5120), .S1(n3929), 
        .Y(n3797) );
  MX4XL U5618 ( .A(\ImageBuffer[52][1] ), .B(\ImageBuffer[53][1] ), .C(
        \ImageBuffer[54][1] ), .D(\ImageBuffer[55][1] ), .S0(n3939), .S1(n3925), .Y(n3782) );
  MX4XL U5619 ( .A(\ImageBuffer[36][1] ), .B(\ImageBuffer[37][1] ), .C(
        \ImageBuffer[38][1] ), .D(\ImageBuffer[39][1] ), .S0(n3939), .S1(n3499), .Y(n3787) );
  MX4XL U5620 ( .A(\ImageBuffer[8][1] ), .B(\ImageBuffer[9][1] ), .C(
        \ImageBuffer[10][1] ), .D(\ImageBuffer[11][1] ), .S0(n5120), .S1(n3480), .Y(n3796) );
  MX4XL U5621 ( .A(\ImageBuffer[40][1] ), .B(\ImageBuffer[41][1] ), .C(
        \ImageBuffer[42][1] ), .D(\ImageBuffer[43][1] ), .S0(n3939), .S1(n3926), .Y(n3786) );
  MXI2XL U5622 ( .A(\ImageBuffer[63][4] ), .B(n4986), .S0(n5411), .Y(n6387) );
  MXI2XL U5623 ( .A(\ImageBuffer[63][1] ), .B(n5025), .S0(n5411), .Y(n6979) );
  MXI2XL U5624 ( .A(\ImageBuffer[63][5] ), .B(n4974), .S0(n5411), .Y(n6189) );
  MXI2XL U5625 ( .A(\ImageBuffer[63][6] ), .B(n4960), .S0(n5411), .Y(n5993) );
  MXI2XL U5626 ( .A(\ImageBuffer[63][7] ), .B(n4949), .S0(n5411), .Y(n5409) );
  MXI2XL U5627 ( .A(\ImageBuffer[63][3] ), .B(n5000), .S0(n5411), .Y(n6585) );
  MXI2XL U5628 ( .A(\ImageBuffer[8][0] ), .B(n5039), .S0(n4934), .Y(n7904) );
  MXI2XL U5629 ( .A(\ImageBuffer[9][0] ), .B(n5040), .S0(n4933), .Y(n7893) );
  MXI2XL U5630 ( .A(\ImageBuffer[11][0] ), .B(n5039), .S0(n4931), .Y(n7870) );
  MXI2XL U5631 ( .A(\ImageBuffer[36][0] ), .B(n5038), .S0(n4903), .Y(n7559) );
  MXI2XL U5632 ( .A(\ImageBuffer[38][0] ), .B(n5038), .S0(n4901), .Y(n7536) );
  MXI2XL U5633 ( .A(\ImageBuffer[41][0] ), .B(n5038), .S0(n4897), .Y(n7490) );
  MXI2XL U5634 ( .A(\ImageBuffer[43][0] ), .B(n5038), .S0(n4895), .Y(n7467) );
  MXI2XL U5635 ( .A(\ImageBuffer[44][0] ), .B(n5038), .S0(n4894), .Y(n7456) );
  MXI2XL U5636 ( .A(\ImageBuffer[46][0] ), .B(n5038), .S0(n4892), .Y(n7433) );
  MXI2XL U5637 ( .A(\ImageBuffer[2][0] ), .B(n5038), .S0(n4940), .Y(n7988) );
  MXI2XL U5638 ( .A(\ImageBuffer[40][0] ), .B(n5038), .S0(n4898), .Y(n7501) );
  MXI2XL U5639 ( .A(\ImageBuffer[48][0] ), .B(n5039), .S0(n4889), .Y(n7401) );
  MXI2XL U5640 ( .A(\ImageBuffer[49][0] ), .B(n5039), .S0(n4888), .Y(n7390) );
  MXI2XL U5641 ( .A(\ImageBuffer[51][0] ), .B(n5039), .S0(n4886), .Y(n7367) );
  MXI2XL U5642 ( .A(\ImageBuffer[52][0] ), .B(n5039), .S0(n4885), .Y(n7356) );
  MXI2XL U5643 ( .A(\ImageBuffer[54][0] ), .B(n5039), .S0(n4883), .Y(n7333) );
  MXI2XL U5644 ( .A(\ImageBuffer[30][0] ), .B(n5038), .S0(n4910), .Y(n7636) );
  MXI2XL U5645 ( .A(\ImageBuffer[33][0] ), .B(n5039), .S0(n4906), .Y(n7593) );
  MXI2XL U5646 ( .A(\ImageBuffer[35][0] ), .B(n5038), .S0(n4904), .Y(n7570) );
  MXI2XL U5647 ( .A(\ImageBuffer[24][0] ), .B(n5039), .S0(n4916), .Y(n7704) );
  MXI2XL U5648 ( .A(\ImageBuffer[25][0] ), .B(n5038), .S0(n4915), .Y(n7693) );
  MXI2XL U5649 ( .A(\ImageBuffer[27][0] ), .B(n5039), .S0(n4913), .Y(n7670) );
  MXI2XL U5650 ( .A(\ImageBuffer[28][0] ), .B(n5040), .S0(n4912), .Y(n7659) );
  MXI2XL U5651 ( .A(\ImageBuffer[60][4] ), .B(n4986), .S0(n4876), .Y(n6401) );
  MXI2XL U5652 ( .A(\ImageBuffer[62][4] ), .B(n4986), .S0(n4874), .Y(n6395) );
  MXI2XL U5653 ( .A(\ImageBuffer[61][1] ), .B(n5025), .S0(n4875), .Y(n6990) );
  MXI2XL U5654 ( .A(\ImageBuffer[60][1] ), .B(n5025), .S0(n4876), .Y(n6993) );
  MXI2XL U5655 ( .A(\ImageBuffer[62][1] ), .B(n5025), .S0(n4874), .Y(n6987) );
  MXI2XL U5656 ( .A(\ImageBuffer[61][5] ), .B(n4975), .S0(n4875), .Y(n6200) );
  MXI2XL U5657 ( .A(\ImageBuffer[60][5] ), .B(n4974), .S0(n4876), .Y(n6203) );
  MXI2XL U5658 ( .A(\ImageBuffer[60][6] ), .B(n4961), .S0(n4876), .Y(n6005) );
  MXI2XL U5659 ( .A(\ImageBuffer[60][7] ), .B(n4949), .S0(n4876), .Y(n5440) );
  MXI2XL U5660 ( .A(\ImageBuffer[62][5] ), .B(n4975), .S0(n4874), .Y(n6197) );
  MXI2XL U5661 ( .A(\ImageBuffer[62][6] ), .B(n4961), .S0(n4874), .Y(n5999) );
  MXI2XL U5662 ( .A(\ImageBuffer[62][7] ), .B(n4950), .S0(n4874), .Y(n5422) );
  MXI2XL U5663 ( .A(\ImageBuffer[61][3] ), .B(n4998), .S0(n4875), .Y(n6595) );
  MXI2XL U5664 ( .A(\ImageBuffer[60][3] ), .B(n5000), .S0(n4876), .Y(n6598) );
  MXI2XL U5665 ( .A(\ImageBuffer[62][3] ), .B(n4998), .S0(n4874), .Y(n6592) );
  MX4XL U5666 ( .A(\ImageBuffer[12][1] ), .B(\ImageBuffer[13][1] ), .C(
        \ImageBuffer[14][1] ), .D(\ImageBuffer[15][1] ), .S0(n4300), .S1(n4306), .Y(n4172) );
  MX4XL U5667 ( .A(\ImageBuffer[4][1] ), .B(\ImageBuffer[5][1] ), .C(
        \ImageBuffer[6][1] ), .D(\ImageBuffer[7][1] ), .S0(n4300), .S1(n4305), 
        .Y(n4174) );
  MX4XL U5668 ( .A(\ImageBuffer[8][1] ), .B(\ImageBuffer[9][1] ), .C(
        \ImageBuffer[10][1] ), .D(\ImageBuffer[11][1] ), .S0(n4300), .S1(n4313), .Y(n4173) );
  MX4XL U5669 ( .A(\ImageBuffer[12][1] ), .B(\ImageBuffer[13][1] ), .C(
        \ImageBuffer[14][1] ), .D(\ImageBuffer[15][1] ), .S0(n4115), .S1(n5116), .Y(n3983) );
  MX4XL U5670 ( .A(n4011), .B(n4009), .C(n4010), .D(n4008), .S0(n4108), .S1(
        n4135), .Y(n4012) );
  MX4XL U5671 ( .A(\ImageBuffer[56][3] ), .B(\ImageBuffer[57][3] ), .C(
        \ImageBuffer[58][3] ), .D(\ImageBuffer[59][3] ), .S0(n3735), .S1(n4133), .Y(n4009) );
  MX4XL U5672 ( .A(\ImageBuffer[60][3] ), .B(\ImageBuffer[61][3] ), .C(
        \ImageBuffer[62][3] ), .D(\ImageBuffer[63][3] ), .S0(n3735), .S1(n3751), .Y(n4008) );
  MX4XL U5673 ( .A(n3883), .B(n3881), .C(n3882), .D(n3880), .S0(n3933), .S1(
        n3409), .Y(n3884) );
  MX4XL U5674 ( .A(\ImageBuffer[60][3] ), .B(\ImageBuffer[61][3] ), .C(
        \ImageBuffer[62][3] ), .D(\ImageBuffer[63][3] ), .S0(n3939), .S1(n5123), .Y(n3820) );
  MX4XL U5675 ( .A(\ImageBuffer[12][1] ), .B(\ImageBuffer[13][1] ), .C(
        \ImageBuffer[14][1] ), .D(\ImageBuffer[15][1] ), .S0(n3735), .S1(n3755), .Y(n3608) );
  MX4XL U5676 ( .A(\ImageBuffer[44][1] ), .B(\ImageBuffer[45][1] ), .C(
        \ImageBuffer[46][1] ), .D(\ImageBuffer[47][1] ), .S0(n3740), .S1(n3754), .Y(n3598) );
  MX4XL U5677 ( .A(\ImageBuffer[60][3] ), .B(\ImageBuffer[61][3] ), .C(
        \ImageBuffer[62][3] ), .D(\ImageBuffer[63][3] ), .S0(n3506), .S1(n3482), .Y(n4539) );
  MX4XL U5678 ( .A(\ImageBuffer[60][5] ), .B(\ImageBuffer[61][5] ), .C(
        \ImageBuffer[62][5] ), .D(\ImageBuffer[63][5] ), .S0(n3935), .S1(n3932), .Y(n3860) );
  MX4XL U5679 ( .A(\ImageBuffer[44][5] ), .B(\ImageBuffer[45][5] ), .C(
        \ImageBuffer[46][5] ), .D(\ImageBuffer[47][5] ), .S0(n3935), .S1(n3921), .Y(n3865) );
  MX4XL U5680 ( .A(\ImageBuffer[28][1] ), .B(\ImageBuffer[29][1] ), .C(
        \ImageBuffer[30][1] ), .D(\ImageBuffer[31][1] ), .S0(n4300), .S1(n4317), .Y(n4167) );
  MX4XL U5681 ( .A(\ImageBuffer[0][1] ), .B(\ImageBuffer[1][1] ), .C(
        \ImageBuffer[2][1] ), .D(\ImageBuffer[3][1] ), .S0(n4115), .S1(n3749), 
        .Y(n3986) );
  MX4XL U5682 ( .A(\ImageBuffer[0][3] ), .B(\ImageBuffer[1][3] ), .C(
        \ImageBuffer[2][3] ), .D(\ImageBuffer[3][3] ), .S0(n4119), .S1(n3750), 
        .Y(n4026) );
  MX4XL U5683 ( .A(\ImageBuffer[16][0] ), .B(\ImageBuffer[17][0] ), .C(
        \ImageBuffer[18][0] ), .D(\ImageBuffer[19][0] ), .S0(n3740), .S1(n4129), .Y(n3586) );
  MX4XL U5684 ( .A(\ImageBuffer[0][3] ), .B(\ImageBuffer[1][3] ), .C(
        \ImageBuffer[2][3] ), .D(\ImageBuffer[3][3] ), .S0(n3506), .S1(n3484), 
        .Y(n4557) );
  MX4XL U5685 ( .A(\ImageBuffer[0][3] ), .B(\ImageBuffer[1][3] ), .C(
        \ImageBuffer[2][3] ), .D(\ImageBuffer[3][3] ), .S0(n3518), .S1(n3471), 
        .Y(n4397) );
  MX4XL U5686 ( .A(\ImageBuffer[0][3] ), .B(\ImageBuffer[1][3] ), .C(
        \ImageBuffer[2][3] ), .D(\ImageBuffer[3][3] ), .S0(n3486), .S1(n3929), 
        .Y(n3838) );
  MX4XL U5687 ( .A(\ImageBuffer[0][1] ), .B(\ImageBuffer[1][1] ), .C(
        \ImageBuffer[2][1] ), .D(\ImageBuffer[3][1] ), .S0(n3735), .S1(n5116), 
        .Y(n3611) );
  MX4XL U5688 ( .A(\ImageBuffer[32][1] ), .B(\ImageBuffer[33][1] ), .C(
        \ImageBuffer[34][1] ), .D(\ImageBuffer[35][1] ), .S0(n3740), .S1(n3748), .Y(n3601) );
  MX4XL U5689 ( .A(\ImageBuffer[16][5] ), .B(\ImageBuffer[17][5] ), .C(
        \ImageBuffer[18][5] ), .D(\ImageBuffer[19][5] ), .S0(n4300), .S1(n3924), .Y(n3873) );
  MX4XL U5690 ( .A(n3878), .B(n3876), .C(n3877), .D(n3875), .S0(n3933), .S1(
        n3409), .Y(n3879) );
  MX4XL U5691 ( .A(\ImageBuffer[8][5] ), .B(\ImageBuffer[9][5] ), .C(
        \ImageBuffer[10][5] ), .D(\ImageBuffer[11][5] ), .S0(n4300), .S1(n3480), .Y(n3876) );
  MX4XL U5692 ( .A(\ImageBuffer[0][5] ), .B(\ImageBuffer[1][5] ), .C(
        \ImageBuffer[2][5] ), .D(\ImageBuffer[3][5] ), .S0(n4300), .S1(n3340), 
        .Y(n3878) );
  MX4XL U5693 ( .A(\ImageBuffer[48][5] ), .B(\ImageBuffer[49][5] ), .C(
        \ImageBuffer[50][5] ), .D(\ImageBuffer[51][5] ), .S0(n3935), .S1(n3921), .Y(n3863) );
  MX4XL U5694 ( .A(\ImageBuffer[32][5] ), .B(\ImageBuffer[33][5] ), .C(
        \ImageBuffer[34][5] ), .D(\ImageBuffer[35][5] ), .S0(n3935), .S1(n3923), .Y(n3868) );
  MX4XL U5695 ( .A(\ImageBuffer[16][7] ), .B(\ImageBuffer[17][7] ), .C(
        \ImageBuffer[18][7] ), .D(\ImageBuffer[19][7] ), .S0(n3938), .S1(n3921), .Y(n3913) );
  MX4XL U5696 ( .A(\ImageBuffer[16][1] ), .B(\ImageBuffer[17][1] ), .C(
        \ImageBuffer[18][1] ), .D(\ImageBuffer[19][1] ), .S0(n4300), .S1(n4307), .Y(n4170) );
  MX4XL U5697 ( .A(\ImageBuffer[0][1] ), .B(\ImageBuffer[1][1] ), .C(
        \ImageBuffer[2][1] ), .D(\ImageBuffer[3][1] ), .S0(n4300), .S1(n4306), 
        .Y(n4175) );
  MX4XL U5698 ( .A(\ImageBuffer[32][1] ), .B(\ImageBuffer[33][1] ), .C(
        \ImageBuffer[34][1] ), .D(\ImageBuffer[35][1] ), .S0(n3939), .S1(n5113), .Y(n4165) );
  MX4XL U5699 ( .A(\ImageBuffer[16][1] ), .B(\ImageBuffer[17][1] ), .C(
        \ImageBuffer[18][1] ), .D(\ImageBuffer[19][1] ), .S0(n4115), .S1(n3749), .Y(n3981) );
  MX4XL U5700 ( .A(\ImageBuffer[24][1] ), .B(\ImageBuffer[25][1] ), .C(
        \ImageBuffer[26][1] ), .D(\ImageBuffer[27][1] ), .S0(n4115), .S1(n3748), .Y(n3979) );
  MX4XL U5701 ( .A(\ImageBuffer[4][1] ), .B(\ImageBuffer[5][1] ), .C(
        \ImageBuffer[6][1] ), .D(\ImageBuffer[7][1] ), .S0(n4115), .S1(n4127), 
        .Y(n3985) );
  MX4XL U5702 ( .A(n4021), .B(n4019), .C(n4020), .D(n4018), .S0(n4108), .S1(
        n4135), .Y(n4022) );
  MX4XL U5703 ( .A(n3893), .B(n3891), .C(n3892), .D(n3890), .S0(n3933), .S1(
        n3409), .Y(n3894) );
  MX4XL U5704 ( .A(\ImageBuffer[16][1] ), .B(\ImageBuffer[17][1] ), .C(
        \ImageBuffer[18][1] ), .D(\ImageBuffer[19][1] ), .S0(n3736), .S1(n4126), .Y(n3606) );
  MX4XL U5705 ( .A(\ImageBuffer[24][1] ), .B(\ImageBuffer[25][1] ), .C(
        \ImageBuffer[26][1] ), .D(\ImageBuffer[27][1] ), .S0(n3736), .S1(n4127), .Y(n3604) );
  MX4XL U5706 ( .A(\ImageBuffer[28][1] ), .B(\ImageBuffer[29][1] ), .C(
        \ImageBuffer[30][1] ), .D(\ImageBuffer[31][1] ), .S0(n3736), .S1(n3747), .Y(n3603) );
  MX4XL U5707 ( .A(\ImageBuffer[4][1] ), .B(\ImageBuffer[5][1] ), .C(
        \ImageBuffer[6][1] ), .D(\ImageBuffer[7][1] ), .S0(n3735), .S1(n3749), 
        .Y(n3610) );
  MX4XL U5708 ( .A(\ImageBuffer[36][1] ), .B(\ImageBuffer[37][1] ), .C(
        \ImageBuffer[38][1] ), .D(\ImageBuffer[39][1] ), .S0(n3740), .S1(n3750), .Y(n3600) );
  MX4XL U5709 ( .A(n3873), .B(n3871), .C(n3872), .D(n3870), .S0(n3933), .S1(
        n3409), .Y(n3874) );
  MX4XL U5710 ( .A(\ImageBuffer[28][5] ), .B(\ImageBuffer[29][5] ), .C(
        \ImageBuffer[30][5] ), .D(\ImageBuffer[31][5] ), .S0(n3935), .S1(n3924), .Y(n3870) );
  MX4XL U5711 ( .A(\ImageBuffer[24][5] ), .B(\ImageBuffer[25][5] ), .C(
        \ImageBuffer[26][5] ), .D(\ImageBuffer[27][5] ), .S0(n4300), .S1(n3921), .Y(n3871) );
  MX4XL U5712 ( .A(\ImageBuffer[52][5] ), .B(\ImageBuffer[53][5] ), .C(
        \ImageBuffer[54][5] ), .D(\ImageBuffer[55][5] ), .S0(n3935), .S1(n3926), .Y(n3862) );
  MX4XL U5713 ( .A(\ImageBuffer[36][5] ), .B(\ImageBuffer[37][5] ), .C(
        \ImageBuffer[38][5] ), .D(\ImageBuffer[39][5] ), .S0(n3935), .S1(n5123), .Y(n3867) );
  MX4XL U5714 ( .A(\ImageBuffer[20][1] ), .B(\ImageBuffer[21][1] ), .C(
        \ImageBuffer[22][1] ), .D(\ImageBuffer[23][1] ), .S0(n4115), .S1(n3752), .Y(n3980) );
  MX4XL U5715 ( .A(\ImageBuffer[52][1] ), .B(\ImageBuffer[53][1] ), .C(
        \ImageBuffer[54][1] ), .D(\ImageBuffer[55][1] ), .S0(n3740), .S1(n4128), .Y(n3595) );
  MX4XL U5716 ( .A(\ImageBuffer[20][1] ), .B(\ImageBuffer[21][1] ), .C(
        \ImageBuffer[22][1] ), .D(\ImageBuffer[23][1] ), .S0(n4300), .S1(n4305), .Y(n4169) );
  MX4XL U5717 ( .A(\ImageBuffer[52][1] ), .B(\ImageBuffer[53][1] ), .C(
        \ImageBuffer[54][1] ), .D(\ImageBuffer[55][1] ), .S0(n3939), .S1(n5113), .Y(n4159) );
  MX4XL U5718 ( .A(\ImageBuffer[8][1] ), .B(\ImageBuffer[9][1] ), .C(
        \ImageBuffer[10][1] ), .D(\ImageBuffer[11][1] ), .S0(n4115), .S1(n3751), .Y(n3984) );
  MX4XL U5719 ( .A(n4016), .B(n4014), .C(n4015), .D(n4013), .S0(n4108), .S1(
        n4135), .Y(n4017) );
  MX4XL U5720 ( .A(\ImageBuffer[56][3] ), .B(\ImageBuffer[57][3] ), .C(
        \ImageBuffer[58][3] ), .D(\ImageBuffer[59][3] ), .S0(n3939), .S1(n3926), .Y(n3821) );
  MX4XL U5721 ( .A(\ImageBuffer[8][1] ), .B(\ImageBuffer[9][1] ), .C(
        \ImageBuffer[10][1] ), .D(\ImageBuffer[11][1] ), .S0(n3735), .S1(n4122), .Y(n3609) );
  MX4XL U5722 ( .A(\ImageBuffer[40][1] ), .B(\ImageBuffer[41][1] ), .C(
        \ImageBuffer[42][1] ), .D(\ImageBuffer[43][1] ), .S0(n3740), .S1(n3757), .Y(n3599) );
  MX4XL U5723 ( .A(\ImageBuffer[56][5] ), .B(\ImageBuffer[57][5] ), .C(
        \ImageBuffer[58][5] ), .D(\ImageBuffer[59][5] ), .S0(n3935), .S1(n3920), .Y(n3861) );
  MX4XL U5724 ( .A(\ImageBuffer[40][5] ), .B(\ImageBuffer[41][5] ), .C(
        \ImageBuffer[42][5] ), .D(\ImageBuffer[43][5] ), .S0(n3935), .S1(n3927), .Y(n3866) );
  MX4XL U5725 ( .A(\ImageBuffer[24][1] ), .B(\ImageBuffer[25][1] ), .C(
        \ImageBuffer[26][1] ), .D(\ImageBuffer[27][1] ), .S0(n4300), .S1(n4303), .Y(n4168) );
  MX4XL U5726 ( .A(\ImageBuffer[40][1] ), .B(\ImageBuffer[41][1] ), .C(
        \ImageBuffer[42][1] ), .D(\ImageBuffer[43][1] ), .S0(n3939), .S1(n4308), .Y(n4163) );
  MX4XL U5727 ( .A(\ImageBuffer[20][1] ), .B(\ImageBuffer[21][1] ), .C(
        \ImageBuffer[22][1] ), .D(\ImageBuffer[23][1] ), .S0(n3516), .S1(n3471), .Y(n4351) );
  MX4X2 U5728 ( .A(n4352), .B(n4350), .C(n4351), .D(n4349), .S0(n3503), .S1(
        n3495), .Y(n4353) );
  MX4XL U5729 ( .A(\ImageBuffer[16][0] ), .B(\ImageBuffer[17][0] ), .C(
        \ImageBuffer[18][0] ), .D(\ImageBuffer[19][0] ), .S0(n3735), .S1(n3749), .Y(n3961) );
  MX4XL U5730 ( .A(\ImageBuffer[52][1] ), .B(\ImageBuffer[53][1] ), .C(
        \ImageBuffer[54][1] ), .D(\ImageBuffer[55][1] ), .S0(n3735), .S1(N2494), .Y(n3970) );
  MX4XL U5731 ( .A(\ImageBuffer[36][1] ), .B(\ImageBuffer[37][1] ), .C(
        \ImageBuffer[38][1] ), .D(\ImageBuffer[39][1] ), .S0(n3735), .S1(n3749), .Y(n3975) );
  MX4X2 U5732 ( .A(n3596), .B(n3594), .C(n3595), .D(n3593), .S0(n3733), .S1(
        n3759), .Y(n3597) );
  MX4XL U5733 ( .A(\ImageBuffer[48][1] ), .B(\ImageBuffer[49][1] ), .C(
        \ImageBuffer[50][1] ), .D(\ImageBuffer[51][1] ), .S0(n3740), .S1(n4122), .Y(n3596) );
  MX4XL U5734 ( .A(\ImageBuffer[56][1] ), .B(\ImageBuffer[57][1] ), .C(
        \ImageBuffer[58][1] ), .D(\ImageBuffer[59][1] ), .S0(n3740), .S1(n3749), .Y(n3594) );
  MX4XL U5735 ( .A(\ImageBuffer[60][1] ), .B(\ImageBuffer[61][1] ), .C(
        \ImageBuffer[62][1] ), .D(\ImageBuffer[63][1] ), .S0(n3740), .S1(n4132), .Y(n3593) );
  MX4X2 U5736 ( .A(n3586), .B(n3584), .C(n3585), .D(n3583), .S0(n3733), .S1(
        n3759), .Y(n3587) );
  MX4XL U5737 ( .A(n3903), .B(n3901), .C(n3902), .D(n3900), .S0(n3933), .S1(
        n3409), .Y(n3904) );
  MX4XL U5738 ( .A(\ImageBuffer[60][7] ), .B(\ImageBuffer[61][7] ), .C(
        \ImageBuffer[62][7] ), .D(\ImageBuffer[63][7] ), .S0(n3939), .S1(n3925), .Y(n3900) );
  MX4XL U5739 ( .A(\ImageBuffer[52][7] ), .B(\ImageBuffer[53][7] ), .C(
        \ImageBuffer[54][7] ), .D(\ImageBuffer[55][7] ), .S0(n3939), .S1(n3921), .Y(n3902) );
  MX4XL U5740 ( .A(\ImageBuffer[56][7] ), .B(\ImageBuffer[57][7] ), .C(
        \ImageBuffer[58][7] ), .D(\ImageBuffer[59][7] ), .S0(n3935), .S1(n3499), .Y(n3901) );
  MX4XL U5741 ( .A(\ImageBuffer[60][3] ), .B(\ImageBuffer[61][3] ), .C(
        \ImageBuffer[62][3] ), .D(\ImageBuffer[63][3] ), .S0(n3938), .S1(n4310), .Y(n4197) );
  MX4XL U5742 ( .A(\ImageBuffer[56][3] ), .B(\ImageBuffer[57][3] ), .C(
        \ImageBuffer[58][3] ), .D(\ImageBuffer[59][3] ), .S0(n3938), .S1(n4313), .Y(n4198) );
  MX4XL U5743 ( .A(n3913), .B(n3911), .C(n3912), .D(n3910), .S0(n3933), .S1(
        n3409), .Y(n3914) );
  MX4XL U5744 ( .A(n4290), .B(n4288), .C(n4289), .D(n4287), .S0(n5108), .S1(
        n3487), .Y(n4291) );
  MX4XL U5745 ( .A(n4255), .B(n4253), .C(n4254), .D(n4252), .S0(n5108), .S1(
        n3487), .Y(n4256) );
  MX4XL U5746 ( .A(\ImageBuffer[12][5] ), .B(\ImageBuffer[13][5] ), .C(
        \ImageBuffer[14][5] ), .D(\ImageBuffer[15][5] ), .S0(n4301), .S1(n4310), .Y(n4252) );
  MX4XL U5747 ( .A(\ImageBuffer[4][5] ), .B(\ImageBuffer[5][5] ), .C(
        \ImageBuffer[6][5] ), .D(\ImageBuffer[7][5] ), .S0(n4301), .S1(n4315), 
        .Y(n4254) );
  MX4XL U5748 ( .A(\ImageBuffer[8][5] ), .B(\ImageBuffer[9][5] ), .C(
        \ImageBuffer[10][5] ), .D(\ImageBuffer[11][5] ), .S0(n4301), .S1(n4310), .Y(n4253) );
  MX4XL U5749 ( .A(n4091), .B(n4089), .C(n4090), .D(n4088), .S0(n4109), .S1(
        n4136), .Y(n4092) );
  MX4XL U5750 ( .A(\ImageBuffer[56][7] ), .B(\ImageBuffer[57][7] ), .C(
        \ImageBuffer[58][7] ), .D(\ImageBuffer[59][7] ), .S0(n4118), .S1(n4123), .Y(n4089) );
  MX4XL U5751 ( .A(\ImageBuffer[60][7] ), .B(\ImageBuffer[61][7] ), .C(
        \ImageBuffer[62][7] ), .D(\ImageBuffer[63][7] ), .S0(n4118), .S1(n4130), .Y(n4088) );
  MX4XL U5752 ( .A(\ImageBuffer[48][5] ), .B(\ImageBuffer[49][5] ), .C(
        \ImageBuffer[50][5] ), .D(\ImageBuffer[51][5] ), .S0(n3743), .S1(n3753), .Y(n4051) );
  MX4XL U5753 ( .A(\ImageBuffer[56][5] ), .B(\ImageBuffer[57][5] ), .C(
        \ImageBuffer[58][5] ), .D(\ImageBuffer[59][5] ), .S0(n3743), .S1(n4128), .Y(n4049) );
  MX4XL U5754 ( .A(\ImageBuffer[60][5] ), .B(\ImageBuffer[61][5] ), .C(
        \ImageBuffer[62][5] ), .D(\ImageBuffer[63][5] ), .S0(n3743), .S1(n4128), .Y(n4048) );
  MX4XL U5755 ( .A(\ImageBuffer[44][5] ), .B(\ImageBuffer[45][5] ), .C(
        \ImageBuffer[46][5] ), .D(\ImageBuffer[47][5] ), .S0(n3743), .S1(n4129), .Y(n4053) );
  MX4XL U5756 ( .A(n3676), .B(n3674), .C(n3675), .D(n3673), .S0(n3734), .S1(
        n3759), .Y(n3677) );
  MX4XL U5757 ( .A(\ImageBuffer[48][5] ), .B(\ImageBuffer[49][5] ), .C(
        \ImageBuffer[50][5] ), .D(\ImageBuffer[51][5] ), .S0(n4116), .S1(n3749), .Y(n3676) );
  MX4XL U5758 ( .A(\ImageBuffer[56][5] ), .B(\ImageBuffer[57][5] ), .C(
        \ImageBuffer[58][5] ), .D(\ImageBuffer[59][5] ), .S0(n4116), .S1(n3754), .Y(n3674) );
  MX4XL U5759 ( .A(\ImageBuffer[60][5] ), .B(\ImageBuffer[61][5] ), .C(
        \ImageBuffer[62][5] ), .D(\ImageBuffer[63][5] ), .S0(n3737), .S1(n4127), .Y(n3673) );
  MX4XL U5760 ( .A(\ImageBuffer[44][5] ), .B(\ImageBuffer[45][5] ), .C(
        \ImageBuffer[46][5] ), .D(\ImageBuffer[47][5] ), .S0(n3498), .S1(n3756), .Y(n3678) );
  MX4XL U5761 ( .A(\ImageBuffer[12][5] ), .B(\ImageBuffer[13][5] ), .C(
        \ImageBuffer[14][5] ), .D(\ImageBuffer[15][5] ), .S0(n3743), .S1(n3747), .Y(n3688) );
  MX4XL U5762 ( .A(\ImageBuffer[60][5] ), .B(\ImageBuffer[61][5] ), .C(
        \ImageBuffer[62][5] ), .D(\ImageBuffer[63][5] ), .S0(n3939), .S1(n4308), .Y(n4237) );
  MX4XL U5763 ( .A(\ImageBuffer[44][5] ), .B(\ImageBuffer[45][5] ), .C(
        \ImageBuffer[46][5] ), .D(\ImageBuffer[47][5] ), .S0(n3939), .S1(n4306), .Y(n4242) );
  MX4XL U5764 ( .A(\ImageBuffer[28][5] ), .B(\ImageBuffer[29][5] ), .C(
        \ImageBuffer[30][5] ), .D(\ImageBuffer[31][5] ), .S0(n4298), .S1(n4314), .Y(n4247) );
  MX4XL U5765 ( .A(\ImageBuffer[60][7] ), .B(\ImageBuffer[61][7] ), .C(
        \ImageBuffer[62][7] ), .D(\ImageBuffer[63][7] ), .S0(n4301), .S1(n4313), .Y(n4277) );
  MX4XL U5766 ( .A(\ImageBuffer[32][5] ), .B(\ImageBuffer[33][5] ), .C(
        \ImageBuffer[34][5] ), .D(\ImageBuffer[35][5] ), .S0(n3743), .S1(n4130), .Y(n4056) );
  MX4XL U5767 ( .A(\ImageBuffer[32][5] ), .B(\ImageBuffer[33][5] ), .C(
        \ImageBuffer[34][5] ), .D(\ImageBuffer[35][5] ), .S0(n4112), .S1(n4125), .Y(n3681) );
  MX4XL U5768 ( .A(\ImageBuffer[0][5] ), .B(\ImageBuffer[1][5] ), .C(
        \ImageBuffer[2][5] ), .D(\ImageBuffer[3][5] ), .S0(n3743), .S1(n4128), 
        .Y(n3691) );
  MX4XL U5769 ( .A(\ImageBuffer[0][5] ), .B(\ImageBuffer[1][5] ), .C(
        \ImageBuffer[2][5] ), .D(\ImageBuffer[3][5] ), .S0(n4301), .S1(n4317), 
        .Y(n4255) );
  MX4XL U5770 ( .A(\ImageBuffer[48][5] ), .B(\ImageBuffer[49][5] ), .C(
        \ImageBuffer[50][5] ), .D(\ImageBuffer[51][5] ), .S0(n4298), .S1(n4314), .Y(n4240) );
  MX4XL U5771 ( .A(\ImageBuffer[32][5] ), .B(\ImageBuffer[33][5] ), .C(
        \ImageBuffer[34][5] ), .D(\ImageBuffer[35][5] ), .S0(n4298), .S1(n4304), .Y(n4245) );
  MX4XL U5772 ( .A(\ImageBuffer[16][5] ), .B(\ImageBuffer[17][5] ), .C(
        \ImageBuffer[18][5] ), .D(\ImageBuffer[19][5] ), .S0(n4301), .S1(n4304), .Y(n4250) );
  MX4XL U5773 ( .A(n4101), .B(n4099), .C(n4100), .D(n4098), .S0(n4109), .S1(
        n4136), .Y(n4102) );
  MX4XL U5774 ( .A(\ImageBuffer[28][5] ), .B(\ImageBuffer[29][5] ), .C(
        \ImageBuffer[30][5] ), .D(\ImageBuffer[31][5] ), .S0(n3743), .S1(n4133), .Y(n4058) );
  MX4XL U5775 ( .A(\ImageBuffer[36][5] ), .B(\ImageBuffer[37][5] ), .C(
        \ImageBuffer[38][5] ), .D(\ImageBuffer[39][5] ), .S0(n3743), .S1(N2494), .Y(n4055) );
  MX4XL U5776 ( .A(n3726), .B(n3724), .C(n3725), .D(n3723), .S0(n3733), .S1(
        n3759), .Y(n3727) );
  MX4XL U5777 ( .A(\ImageBuffer[28][5] ), .B(\ImageBuffer[29][5] ), .C(
        \ImageBuffer[30][5] ), .D(\ImageBuffer[31][5] ), .S0(n4112), .S1(n4124), .Y(n3683) );
  MX4XL U5778 ( .A(\ImageBuffer[36][5] ), .B(\ImageBuffer[37][5] ), .C(
        \ImageBuffer[38][5] ), .D(\ImageBuffer[39][5] ), .S0(n3498), .S1(n5116), .Y(n3680) );
  MX4XL U5779 ( .A(\ImageBuffer[52][5] ), .B(\ImageBuffer[53][5] ), .C(
        \ImageBuffer[54][5] ), .D(\ImageBuffer[55][5] ), .S0(n3743), .S1(n4131), .Y(n4050) );
  MX4XL U5780 ( .A(\ImageBuffer[52][5] ), .B(\ImageBuffer[53][5] ), .C(
        \ImageBuffer[54][5] ), .D(\ImageBuffer[55][5] ), .S0(n4298), .S1(n4310), .Y(n4239) );
  MX4XL U5781 ( .A(\ImageBuffer[36][5] ), .B(\ImageBuffer[37][5] ), .C(
        \ImageBuffer[38][5] ), .D(\ImageBuffer[39][5] ), .S0(n4298), .S1(n4308), .Y(n4244) );
  MX4XL U5782 ( .A(\ImageBuffer[20][5] ), .B(\ImageBuffer[21][5] ), .C(
        \ImageBuffer[22][5] ), .D(\ImageBuffer[23][5] ), .S0(n4301), .S1(n4315), .Y(n4249) );
  MX4XL U5783 ( .A(\ImageBuffer[52][5] ), .B(\ImageBuffer[53][5] ), .C(
        \ImageBuffer[54][5] ), .D(\ImageBuffer[55][5] ), .S0(n4116), .S1(n4131), .Y(n3675) );
  MX4XL U5784 ( .A(\ImageBuffer[52][7] ), .B(\ImageBuffer[53][7] ), .C(
        \ImageBuffer[54][7] ), .D(\ImageBuffer[55][7] ), .S0(n4118), .S1(n3751), .Y(n4090) );
  MX4XL U5785 ( .A(\ImageBuffer[52][7] ), .B(\ImageBuffer[53][7] ), .C(
        \ImageBuffer[54][7] ), .D(\ImageBuffer[55][7] ), .S0(n4301), .S1(n4313), .Y(n4279) );
  MX4XL U5786 ( .A(\ImageBuffer[52][7] ), .B(\ImageBuffer[53][7] ), .C(
        \ImageBuffer[54][7] ), .D(\ImageBuffer[55][7] ), .S0(n3488), .S1(n4133), .Y(n3715) );
  MX4XL U5787 ( .A(n4096), .B(n4094), .C(n4095), .D(n4093), .S0(n4109), .S1(
        n4136), .Y(n4097) );
  MX4XL U5788 ( .A(\ImageBuffer[40][5] ), .B(\ImageBuffer[41][5] ), .C(
        \ImageBuffer[42][5] ), .D(\ImageBuffer[43][5] ), .S0(n3743), .S1(n3755), .Y(n4054) );
  MX4XL U5789 ( .A(\ImageBuffer[40][5] ), .B(\ImageBuffer[41][5] ), .C(
        \ImageBuffer[42][5] ), .D(\ImageBuffer[43][5] ), .S0(n3737), .S1(n4134), .Y(n3679) );
  MX4XL U5790 ( .A(\ImageBuffer[8][5] ), .B(\ImageBuffer[9][5] ), .C(
        \ImageBuffer[10][5] ), .D(\ImageBuffer[11][5] ), .S0(n3743), .S1(N2494), .Y(n3689) );
  MX4XL U5791 ( .A(\ImageBuffer[56][5] ), .B(\ImageBuffer[57][5] ), .C(
        \ImageBuffer[58][5] ), .D(\ImageBuffer[59][5] ), .S0(n4298), .S1(n4304), .Y(n4238) );
  MX4XL U5792 ( .A(\ImageBuffer[40][5] ), .B(\ImageBuffer[41][5] ), .C(
        \ImageBuffer[42][5] ), .D(\ImageBuffer[43][5] ), .S0(n4298), .S1(n5113), .Y(n4243) );
  MX4XL U5793 ( .A(\ImageBuffer[24][5] ), .B(\ImageBuffer[25][5] ), .C(
        \ImageBuffer[26][5] ), .D(\ImageBuffer[27][5] ), .S0(n4301), .S1(n4303), .Y(n4248) );
  MX4XL U5794 ( .A(\ImageBuffer[56][7] ), .B(\ImageBuffer[57][7] ), .C(
        \ImageBuffer[58][7] ), .D(\ImageBuffer[59][7] ), .S0(n4297), .S1(n4309), .Y(n4278) );
  CLKBUFX2 U5795 ( .A(N2486), .Y(n4946) );
  NAND2X4 U5796 ( .A(n3477), .B(cmd[3]), .Y(n8028) );
  NAND2X4 U5797 ( .A(n3475), .B(cmd[3]), .Y(n8030) );
  NAND2XL U5798 ( .A(cmd[0]), .B(n8021), .Y(n8015) );
  MX4XL U5799 ( .A(\ImageBuffer[12][0] ), .B(\ImageBuffer[13][0] ), .C(
        \ImageBuffer[14][0] ), .D(\ImageBuffer[15][0] ), .S0(n4803), .S1(n4811), .Y(n4657) );
  MX4XL U5800 ( .A(\ImageBuffer[60][1] ), .B(\ImageBuffer[61][1] ), .C(
        \ImageBuffer[62][1] ), .D(\ImageBuffer[63][1] ), .S0(n4803), .S1(n4811), .Y(n4662) );
  MX4XL U5801 ( .A(\ImageBuffer[44][1] ), .B(\ImageBuffer[45][1] ), .C(
        \ImageBuffer[46][1] ), .D(\ImageBuffer[47][1] ), .S0(n4803), .S1(n4811), .Y(n4667) );
  MX4XL U5802 ( .A(\ImageBuffer[12][1] ), .B(\ImageBuffer[13][1] ), .C(
        \ImageBuffer[14][1] ), .D(\ImageBuffer[15][1] ), .S0(n4804), .S1(n4812), .Y(n4677) );
  MX4XL U5803 ( .A(\ImageBuffer[60][2] ), .B(\ImageBuffer[61][2] ), .C(
        \ImageBuffer[62][2] ), .D(\ImageBuffer[63][2] ), .S0(n4804), .S1(n4812), .Y(n4682) );
  MX4XL U5804 ( .A(\ImageBuffer[44][2] ), .B(\ImageBuffer[45][2] ), .C(
        \ImageBuffer[46][2] ), .D(\ImageBuffer[47][2] ), .S0(n4804), .S1(n4812), .Y(n4687) );
  MX4XL U5805 ( .A(\ImageBuffer[12][2] ), .B(\ImageBuffer[13][2] ), .C(
        \ImageBuffer[14][2] ), .D(\ImageBuffer[15][2] ), .S0(n4805), .S1(n4813), .Y(n4697) );
  MX4XL U5806 ( .A(\ImageBuffer[60][3] ), .B(\ImageBuffer[61][3] ), .C(
        \ImageBuffer[62][3] ), .D(\ImageBuffer[63][3] ), .S0(n4805), .S1(n4813), .Y(n4702) );
  MX4XL U5807 ( .A(\ImageBuffer[44][3] ), .B(\ImageBuffer[45][3] ), .C(
        \ImageBuffer[46][3] ), .D(\ImageBuffer[47][3] ), .S0(n4806), .S1(n4814), .Y(n4707) );
  MX4XL U5808 ( .A(\ImageBuffer[12][3] ), .B(\ImageBuffer[13][3] ), .C(
        \ImageBuffer[14][3] ), .D(\ImageBuffer[15][3] ), .S0(n4806), .S1(n4814), .Y(n4717) );
  MX4XL U5809 ( .A(\ImageBuffer[60][4] ), .B(\ImageBuffer[61][4] ), .C(
        \ImageBuffer[62][4] ), .D(\ImageBuffer[63][4] ), .S0(n4807), .S1(n4812), .Y(n4722) );
  MX4XL U5810 ( .A(\ImageBuffer[44][4] ), .B(\ImageBuffer[45][4] ), .C(
        \ImageBuffer[46][4] ), .D(\ImageBuffer[47][4] ), .S0(n4807), .S1(n4813), .Y(n4727) );
  MX4XL U5811 ( .A(\ImageBuffer[12][4] ), .B(\ImageBuffer[13][4] ), .C(
        \ImageBuffer[14][4] ), .D(\ImageBuffer[15][4] ), .S0(n4806), .S1(n4815), .Y(n4737) );
  MX4XL U5812 ( .A(\ImageBuffer[60][5] ), .B(\ImageBuffer[61][5] ), .C(
        \ImageBuffer[62][5] ), .D(\ImageBuffer[63][5] ), .S0(n4803), .S1(n4815), .Y(n4742) );
  MX4XL U5813 ( .A(\ImageBuffer[44][5] ), .B(\ImageBuffer[45][5] ), .C(
        \ImageBuffer[46][5] ), .D(\ImageBuffer[47][5] ), .S0(n4805), .S1(n4815), .Y(n4747) );
  MX4XL U5814 ( .A(\ImageBuffer[12][5] ), .B(\ImageBuffer[13][5] ), .C(
        \ImageBuffer[14][5] ), .D(\ImageBuffer[15][5] ), .S0(n4804), .S1(n4816), .Y(n4757) );
  MX4XL U5815 ( .A(\ImageBuffer[60][6] ), .B(\ImageBuffer[61][6] ), .C(
        \ImageBuffer[62][6] ), .D(\ImageBuffer[63][6] ), .S0(n4807), .S1(n4816), .Y(n4762) );
  MX4XL U5816 ( .A(\ImageBuffer[44][6] ), .B(\ImageBuffer[45][6] ), .C(
        \ImageBuffer[46][6] ), .D(\ImageBuffer[47][6] ), .S0(n4804), .S1(n4816), .Y(n4767) );
  MX4XL U5817 ( .A(\ImageBuffer[12][6] ), .B(\ImageBuffer[13][6] ), .C(
        \ImageBuffer[14][6] ), .D(\ImageBuffer[15][6] ), .S0(n4808), .S1(n4817), .Y(n4777) );
  MX4XL U5818 ( .A(\ImageBuffer[60][7] ), .B(\ImageBuffer[61][7] ), .C(
        \ImageBuffer[62][7] ), .D(\ImageBuffer[63][7] ), .S0(n4808), .S1(n4817), .Y(n4782) );
  MX4XL U5819 ( .A(\ImageBuffer[44][7] ), .B(\ImageBuffer[45][7] ), .C(
        \ImageBuffer[46][7] ), .D(\ImageBuffer[47][7] ), .S0(n4809), .S1(n4816), .Y(n4787) );
  MX4XL U5820 ( .A(\ImageBuffer[12][7] ), .B(\ImageBuffer[13][7] ), .C(
        \ImageBuffer[14][7] ), .D(\ImageBuffer[15][7] ), .S0(n4809), .S1(n4811), .Y(n4797) );
  MX4XL U5821 ( .A(\ImageBuffer[16][5] ), .B(\ImageBuffer[17][5] ), .C(
        \ImageBuffer[18][5] ), .D(\ImageBuffer[19][5] ), .S0(n4803), .S1(n4816), .Y(n4755) );
  MX4XL U5822 ( .A(\ImageBuffer[24][5] ), .B(\ImageBuffer[25][5] ), .C(
        \ImageBuffer[26][5] ), .D(\ImageBuffer[27][5] ), .S0(n4805), .S1(n4816), .Y(n4753) );
  MX4XL U5823 ( .A(\ImageBuffer[28][5] ), .B(\ImageBuffer[29][5] ), .C(
        \ImageBuffer[30][5] ), .D(\ImageBuffer[31][5] ), .S0(n4807), .S1(n4815), .Y(n4752) );
  MX4XL U5824 ( .A(\ImageBuffer[16][6] ), .B(\ImageBuffer[17][6] ), .C(
        \ImageBuffer[18][6] ), .D(\ImageBuffer[19][6] ), .S0(n4808), .S1(n4817), .Y(n4775) );
  MX4XL U5825 ( .A(\ImageBuffer[24][6] ), .B(\ImageBuffer[25][6] ), .C(
        \ImageBuffer[26][6] ), .D(\ImageBuffer[27][6] ), .S0(n4808), .S1(n4817), .Y(n4773) );
  MX4XL U5826 ( .A(\ImageBuffer[28][6] ), .B(\ImageBuffer[29][6] ), .C(
        \ImageBuffer[30][6] ), .D(\ImageBuffer[31][6] ), .S0(n4808), .S1(n4817), .Y(n4772) );
  MX4XL U5827 ( .A(\ImageBuffer[16][7] ), .B(\ImageBuffer[17][7] ), .C(
        \ImageBuffer[18][7] ), .D(\ImageBuffer[19][7] ), .S0(n4809), .S1(n4810), .Y(n4795) );
  MX4XL U5828 ( .A(\ImageBuffer[24][7] ), .B(\ImageBuffer[25][7] ), .C(
        \ImageBuffer[26][7] ), .D(\ImageBuffer[27][7] ), .S0(n4809), .S1(n4810), .Y(n4793) );
  MX4XL U5829 ( .A(\ImageBuffer[28][7] ), .B(\ImageBuffer[29][7] ), .C(
        \ImageBuffer[30][7] ), .D(\ImageBuffer[31][7] ), .S0(n4809), .S1(n4817), .Y(n4792) );
  MX4XL U5830 ( .A(\ImageBuffer[16][0] ), .B(\ImageBuffer[17][0] ), .C(
        \ImageBuffer[18][0] ), .D(\ImageBuffer[19][0] ), .S0(n4803), .S1(n4811), .Y(n4655) );
  MX4XL U5831 ( .A(\ImageBuffer[0][0] ), .B(\ImageBuffer[1][0] ), .C(
        \ImageBuffer[2][0] ), .D(\ImageBuffer[3][0] ), .S0(n4803), .S1(n4811), 
        .Y(n4660) );
  MX4XL U5832 ( .A(\ImageBuffer[48][1] ), .B(\ImageBuffer[49][1] ), .C(
        \ImageBuffer[50][1] ), .D(\ImageBuffer[51][1] ), .S0(n4803), .S1(n4811), .Y(n4665) );
  MX4XL U5833 ( .A(\ImageBuffer[32][1] ), .B(\ImageBuffer[33][1] ), .C(
        \ImageBuffer[34][1] ), .D(\ImageBuffer[35][1] ), .S0(n4803), .S1(n4811), .Y(n4670) );
  MX4XL U5834 ( .A(\ImageBuffer[0][1] ), .B(\ImageBuffer[1][1] ), .C(
        \ImageBuffer[2][1] ), .D(\ImageBuffer[3][1] ), .S0(n4804), .S1(n4812), 
        .Y(n4680) );
  MX4XL U5835 ( .A(\ImageBuffer[48][2] ), .B(\ImageBuffer[49][2] ), .C(
        \ImageBuffer[50][2] ), .D(\ImageBuffer[51][2] ), .S0(n4804), .S1(n4812), .Y(n4685) );
  MX4XL U5836 ( .A(\ImageBuffer[32][2] ), .B(\ImageBuffer[33][2] ), .C(
        \ImageBuffer[34][2] ), .D(\ImageBuffer[35][2] ), .S0(n4805), .S1(n4813), .Y(n4690) );
  MX4XL U5837 ( .A(\ImageBuffer[0][2] ), .B(\ImageBuffer[1][2] ), .C(
        \ImageBuffer[2][2] ), .D(\ImageBuffer[3][2] ), .S0(n4805), .S1(n4813), 
        .Y(n4700) );
  MX4XL U5838 ( .A(\ImageBuffer[48][3] ), .B(\ImageBuffer[49][3] ), .C(
        \ImageBuffer[50][3] ), .D(\ImageBuffer[51][3] ), .S0(n4806), .S1(n4814), .Y(n4705) );
  MX4XL U5839 ( .A(\ImageBuffer[32][3] ), .B(\ImageBuffer[33][3] ), .C(
        \ImageBuffer[34][3] ), .D(\ImageBuffer[35][3] ), .S0(n4806), .S1(n4814), .Y(n4710) );
  MX4XL U5840 ( .A(\ImageBuffer[0][3] ), .B(\ImageBuffer[1][3] ), .C(
        \ImageBuffer[2][3] ), .D(\ImageBuffer[3][3] ), .S0(n4807), .S1(n4813), 
        .Y(n4720) );
  MX4XL U5841 ( .A(\ImageBuffer[48][4] ), .B(\ImageBuffer[49][4] ), .C(
        \ImageBuffer[50][4] ), .D(\ImageBuffer[51][4] ), .S0(n4807), .S1(n4814), .Y(n4725) );
  MX4XL U5842 ( .A(\ImageBuffer[32][4] ), .B(\ImageBuffer[33][4] ), .C(
        \ImageBuffer[34][4] ), .D(\ImageBuffer[35][4] ), .S0(n4807), .S1(n4812), .Y(n4730) );
  MX4XL U5843 ( .A(\ImageBuffer[0][4] ), .B(\ImageBuffer[1][4] ), .C(
        \ImageBuffer[2][4] ), .D(\ImageBuffer[3][4] ), .S0(n4809), .S1(n4815), 
        .Y(n4740) );
  MX4XL U5844 ( .A(\ImageBuffer[48][5] ), .B(\ImageBuffer[49][5] ), .C(
        \ImageBuffer[50][5] ), .D(\ImageBuffer[51][5] ), .S0(n4806), .S1(n4815), .Y(n4745) );
  MX4XL U5845 ( .A(\ImageBuffer[32][5] ), .B(\ImageBuffer[33][5] ), .C(
        \ImageBuffer[34][5] ), .D(\ImageBuffer[35][5] ), .S0(n4802), .S1(n4815), .Y(n4750) );
  MX4XL U5846 ( .A(\ImageBuffer[0][5] ), .B(\ImageBuffer[1][5] ), .C(
        \ImageBuffer[2][5] ), .D(\ImageBuffer[3][5] ), .S0(n4805), .S1(n4816), 
        .Y(n4760) );
  MX4XL U5847 ( .A(\ImageBuffer[48][6] ), .B(\ImageBuffer[49][6] ), .C(
        \ImageBuffer[50][6] ), .D(\ImageBuffer[51][6] ), .S0(n4807), .S1(n4816), .Y(n4765) );
  MX4XL U5848 ( .A(\ImageBuffer[32][6] ), .B(\ImageBuffer[33][6] ), .C(
        \ImageBuffer[34][6] ), .D(\ImageBuffer[35][6] ), .S0(n4808), .S1(n4817), .Y(n4770) );
  MX4XL U5849 ( .A(\ImageBuffer[0][6] ), .B(\ImageBuffer[1][6] ), .C(
        \ImageBuffer[2][6] ), .D(\ImageBuffer[3][6] ), .S0(n4808), .S1(n4817), 
        .Y(n4780) );
  MX4XL U5850 ( .A(\ImageBuffer[48][7] ), .B(\ImageBuffer[49][7] ), .C(
        \ImageBuffer[50][7] ), .D(\ImageBuffer[51][7] ), .S0(n4809), .S1(n4810), .Y(n4785) );
  MX4XL U5851 ( .A(\ImageBuffer[32][7] ), .B(\ImageBuffer[33][7] ), .C(
        \ImageBuffer[34][7] ), .D(\ImageBuffer[35][7] ), .S0(n4809), .S1(n4810), .Y(n4790) );
  MX4XL U5852 ( .A(\ImageBuffer[0][7] ), .B(\ImageBuffer[1][7] ), .C(
        \ImageBuffer[2][7] ), .D(\ImageBuffer[3][7] ), .S0(n4809), .S1(n4817), 
        .Y(n4800) );
  MX4XL U5853 ( .A(\ImageBuffer[4][0] ), .B(\ImageBuffer[5][0] ), .C(
        \ImageBuffer[6][0] ), .D(\ImageBuffer[7][0] ), .S0(n4803), .S1(n4811), 
        .Y(n4659) );
  MX4XL U5854 ( .A(\ImageBuffer[20][1] ), .B(\ImageBuffer[21][1] ), .C(
        \ImageBuffer[22][1] ), .D(\ImageBuffer[23][1] ), .S0(n4804), .S1(n4812), .Y(n4674) );
  MX4XL U5855 ( .A(\ImageBuffer[52][1] ), .B(\ImageBuffer[53][1] ), .C(
        \ImageBuffer[54][1] ), .D(\ImageBuffer[55][1] ), .S0(n4803), .S1(n4811), .Y(n4664) );
  MX4XL U5856 ( .A(\ImageBuffer[36][1] ), .B(\ImageBuffer[37][1] ), .C(
        \ImageBuffer[38][1] ), .D(\ImageBuffer[39][1] ), .S0(n4803), .S1(n4811), .Y(n4669) );
  MX4XL U5857 ( .A(\ImageBuffer[4][1] ), .B(\ImageBuffer[5][1] ), .C(
        \ImageBuffer[6][1] ), .D(\ImageBuffer[7][1] ), .S0(n4804), .S1(n4812), 
        .Y(n4679) );
  MX4XL U5858 ( .A(\ImageBuffer[20][2] ), .B(\ImageBuffer[21][2] ), .C(
        \ImageBuffer[22][2] ), .D(\ImageBuffer[23][2] ), .S0(n4805), .S1(n4813), .Y(n4694) );
  MX4XL U5859 ( .A(\ImageBuffer[52][2] ), .B(\ImageBuffer[53][2] ), .C(
        \ImageBuffer[54][2] ), .D(\ImageBuffer[55][2] ), .S0(n4804), .S1(n4812), .Y(n4684) );
  MX4XL U5860 ( .A(\ImageBuffer[36][2] ), .B(\ImageBuffer[37][2] ), .C(
        \ImageBuffer[38][2] ), .D(\ImageBuffer[39][2] ), .S0(n4805), .S1(n4813), .Y(n4689) );
  MX4XL U5861 ( .A(\ImageBuffer[4][2] ), .B(\ImageBuffer[5][2] ), .C(
        \ImageBuffer[6][2] ), .D(\ImageBuffer[7][2] ), .S0(n4805), .S1(n4813), 
        .Y(n4699) );
  MX4XL U5862 ( .A(\ImageBuffer[20][3] ), .B(\ImageBuffer[21][3] ), .C(
        \ImageBuffer[22][3] ), .D(\ImageBuffer[23][3] ), .S0(n4806), .S1(n4814), .Y(n4714) );
  MX4XL U5863 ( .A(\ImageBuffer[52][3] ), .B(\ImageBuffer[53][3] ), .C(
        \ImageBuffer[54][3] ), .D(\ImageBuffer[55][3] ), .S0(n4806), .S1(n4814), .Y(n4704) );
  MX4XL U5864 ( .A(\ImageBuffer[36][3] ), .B(\ImageBuffer[37][3] ), .C(
        \ImageBuffer[38][3] ), .D(\ImageBuffer[39][3] ), .S0(n4806), .S1(n4814), .Y(n4709) );
  MX4XL U5865 ( .A(\ImageBuffer[4][3] ), .B(\ImageBuffer[5][3] ), .C(
        \ImageBuffer[6][3] ), .D(\ImageBuffer[7][3] ), .S0(n4806), .S1(n4814), 
        .Y(n4719) );
  MX4XL U5866 ( .A(\ImageBuffer[20][4] ), .B(\ImageBuffer[21][4] ), .C(
        \ImageBuffer[22][4] ), .D(\ImageBuffer[23][4] ), .S0(n4807), .S1(n4812), .Y(n4734) );
  MX4XL U5867 ( .A(\ImageBuffer[52][4] ), .B(\ImageBuffer[53][4] ), .C(
        \ImageBuffer[54][4] ), .D(\ImageBuffer[55][4] ), .S0(n4807), .S1(n4813), .Y(n4724) );
  MX4XL U5868 ( .A(\ImageBuffer[36][4] ), .B(\ImageBuffer[37][4] ), .C(
        \ImageBuffer[38][4] ), .D(\ImageBuffer[39][4] ), .S0(n4807), .S1(n4812), .Y(n4729) );
  MX4XL U5869 ( .A(\ImageBuffer[4][4] ), .B(\ImageBuffer[5][4] ), .C(
        \ImageBuffer[6][4] ), .D(\ImageBuffer[7][4] ), .S0(n4808), .S1(n4815), 
        .Y(n4739) );
  MX4XL U5870 ( .A(\ImageBuffer[20][5] ), .B(\ImageBuffer[21][5] ), .C(
        \ImageBuffer[22][5] ), .D(\ImageBuffer[23][5] ), .S0(n4805), .S1(n4816), .Y(n4754) );
  MX4XL U5871 ( .A(\ImageBuffer[52][5] ), .B(\ImageBuffer[53][5] ), .C(
        \ImageBuffer[54][5] ), .D(\ImageBuffer[55][5] ), .S0(n4803), .S1(n4815), .Y(n4744) );
  MX4XL U5872 ( .A(\ImageBuffer[36][5] ), .B(\ImageBuffer[37][5] ), .C(
        \ImageBuffer[38][5] ), .D(\ImageBuffer[39][5] ), .S0(n4806), .S1(n4815), .Y(n4749) );
  MX4XL U5873 ( .A(\ImageBuffer[4][5] ), .B(\ImageBuffer[5][5] ), .C(
        \ImageBuffer[6][5] ), .D(\ImageBuffer[7][5] ), .S0(n4808), .S1(n4816), 
        .Y(n4759) );
  MX4XL U5874 ( .A(\ImageBuffer[20][6] ), .B(\ImageBuffer[21][6] ), .C(
        \ImageBuffer[22][6] ), .D(\ImageBuffer[23][6] ), .S0(n4808), .S1(n4817), .Y(n4774) );
  MX4XL U5875 ( .A(\ImageBuffer[52][6] ), .B(\ImageBuffer[53][6] ), .C(
        \ImageBuffer[54][6] ), .D(\ImageBuffer[55][6] ), .S0(n4804), .S1(n4816), .Y(n4764) );
  MX4XL U5876 ( .A(\ImageBuffer[36][6] ), .B(\ImageBuffer[37][6] ), .C(
        \ImageBuffer[38][6] ), .D(\ImageBuffer[39][6] ), .S0(n4808), .S1(n4817), .Y(n4769) );
  MX4XL U5877 ( .A(\ImageBuffer[4][6] ), .B(\ImageBuffer[5][6] ), .C(
        \ImageBuffer[6][6] ), .D(\ImageBuffer[7][6] ), .S0(n4808), .S1(n4817), 
        .Y(n4779) );
  MX4XL U5878 ( .A(\ImageBuffer[20][7] ), .B(\ImageBuffer[21][7] ), .C(
        \ImageBuffer[22][7] ), .D(\ImageBuffer[23][7] ), .S0(n4809), .S1(n4815), .Y(n4794) );
  MX4XL U5879 ( .A(\ImageBuffer[52][7] ), .B(\ImageBuffer[53][7] ), .C(
        \ImageBuffer[54][7] ), .D(\ImageBuffer[55][7] ), .S0(n4808), .S1(n4817), .Y(n4784) );
  MX4XL U5880 ( .A(\ImageBuffer[36][7] ), .B(\ImageBuffer[37][7] ), .C(
        \ImageBuffer[38][7] ), .D(\ImageBuffer[39][7] ), .S0(n4809), .S1(n4810), .Y(n4789) );
  MX4XL U5881 ( .A(\ImageBuffer[4][7] ), .B(\ImageBuffer[5][7] ), .C(
        \ImageBuffer[6][7] ), .D(\ImageBuffer[7][7] ), .S0(n4809), .S1(n4812), 
        .Y(n4799) );
  MX4XL U5882 ( .A(\ImageBuffer[16][1] ), .B(\ImageBuffer[17][1] ), .C(
        \ImageBuffer[18][1] ), .D(\ImageBuffer[19][1] ), .S0(n4804), .S1(n4812), .Y(n4675) );
  MX4XL U5883 ( .A(\ImageBuffer[24][1] ), .B(\ImageBuffer[25][1] ), .C(
        \ImageBuffer[26][1] ), .D(\ImageBuffer[27][1] ), .S0(n4804), .S1(n4812), .Y(n4673) );
  MX4XL U5884 ( .A(\ImageBuffer[28][1] ), .B(\ImageBuffer[29][1] ), .C(
        \ImageBuffer[30][1] ), .D(\ImageBuffer[31][1] ), .S0(n4804), .S1(n4812), .Y(n4672) );
  MX4XL U5885 ( .A(\ImageBuffer[16][2] ), .B(\ImageBuffer[17][2] ), .C(
        \ImageBuffer[18][2] ), .D(\ImageBuffer[19][2] ), .S0(n4805), .S1(n4813), .Y(n4695) );
  MX4XL U5886 ( .A(\ImageBuffer[24][2] ), .B(\ImageBuffer[25][2] ), .C(
        \ImageBuffer[26][2] ), .D(\ImageBuffer[27][2] ), .S0(n4805), .S1(n4813), .Y(n4693) );
  MX4XL U5887 ( .A(\ImageBuffer[28][2] ), .B(\ImageBuffer[29][2] ), .C(
        \ImageBuffer[30][2] ), .D(\ImageBuffer[31][2] ), .S0(n4805), .S1(n4813), .Y(n4692) );
  MX4XL U5888 ( .A(\ImageBuffer[16][3] ), .B(\ImageBuffer[17][3] ), .C(
        \ImageBuffer[18][3] ), .D(\ImageBuffer[19][3] ), .S0(n4806), .S1(n4814), .Y(n4715) );
  MX4XL U5889 ( .A(\ImageBuffer[24][3] ), .B(\ImageBuffer[25][3] ), .C(
        \ImageBuffer[26][3] ), .D(\ImageBuffer[27][3] ), .S0(n4806), .S1(n4814), .Y(n4713) );
  MX4XL U5890 ( .A(\ImageBuffer[28][3] ), .B(\ImageBuffer[29][3] ), .C(
        \ImageBuffer[30][3] ), .D(\ImageBuffer[31][3] ), .S0(n4806), .S1(n4814), .Y(n4712) );
  MX4XL U5891 ( .A(\ImageBuffer[16][4] ), .B(\ImageBuffer[17][4] ), .C(
        \ImageBuffer[18][4] ), .D(\ImageBuffer[19][4] ), .S0(n4807), .S1(n4811), .Y(n4735) );
  MX4XL U5892 ( .A(\ImageBuffer[24][4] ), .B(\ImageBuffer[25][4] ), .C(
        \ImageBuffer[26][4] ), .D(\ImageBuffer[27][4] ), .S0(n4807), .S1(n4813), .Y(n4733) );
  MX4XL U5893 ( .A(\ImageBuffer[28][4] ), .B(\ImageBuffer[29][4] ), .C(
        \ImageBuffer[30][4] ), .D(\ImageBuffer[31][4] ), .S0(n4807), .S1(n4811), .Y(n4732) );
  MX4XL U5894 ( .A(\ImageBuffer[8][0] ), .B(\ImageBuffer[9][0] ), .C(
        \ImageBuffer[10][0] ), .D(\ImageBuffer[11][0] ), .S0(n4803), .S1(n4811), .Y(n4658) );
  MX4XL U5895 ( .A(\ImageBuffer[56][1] ), .B(\ImageBuffer[57][1] ), .C(
        \ImageBuffer[58][1] ), .D(\ImageBuffer[59][1] ), .S0(n4803), .S1(n4811), .Y(n4663) );
  MX4XL U5896 ( .A(\ImageBuffer[40][1] ), .B(\ImageBuffer[41][1] ), .C(
        \ImageBuffer[42][1] ), .D(\ImageBuffer[43][1] ), .S0(n4803), .S1(n4811), .Y(n4668) );
  MX4XL U5897 ( .A(\ImageBuffer[8][1] ), .B(\ImageBuffer[9][1] ), .C(
        \ImageBuffer[10][1] ), .D(\ImageBuffer[11][1] ), .S0(n4804), .S1(n4812), .Y(n4678) );
  MX4XL U5898 ( .A(\ImageBuffer[56][2] ), .B(\ImageBuffer[57][2] ), .C(
        \ImageBuffer[58][2] ), .D(\ImageBuffer[59][2] ), .S0(n4804), .S1(n4812), .Y(n4683) );
  MX4XL U5899 ( .A(\ImageBuffer[40][2] ), .B(\ImageBuffer[41][2] ), .C(
        \ImageBuffer[42][2] ), .D(\ImageBuffer[43][2] ), .S0(n4805), .S1(n4813), .Y(n4688) );
  MX4XL U5900 ( .A(\ImageBuffer[8][2] ), .B(\ImageBuffer[9][2] ), .C(
        \ImageBuffer[10][2] ), .D(\ImageBuffer[11][2] ), .S0(n4805), .S1(n4813), .Y(n4698) );
  MX4XL U5901 ( .A(\ImageBuffer[56][3] ), .B(\ImageBuffer[57][3] ), .C(
        \ImageBuffer[58][3] ), .D(\ImageBuffer[59][3] ), .S0(n4805), .S1(n4813), .Y(n4703) );
  MX4XL U5902 ( .A(\ImageBuffer[40][3] ), .B(\ImageBuffer[41][3] ), .C(
        \ImageBuffer[42][3] ), .D(\ImageBuffer[43][3] ), .S0(n4806), .S1(n4814), .Y(n4708) );
  MX4XL U5903 ( .A(\ImageBuffer[8][3] ), .B(\ImageBuffer[9][3] ), .C(
        \ImageBuffer[10][3] ), .D(\ImageBuffer[11][3] ), .S0(n4806), .S1(n4814), .Y(n4718) );
  MX4XL U5904 ( .A(\ImageBuffer[56][4] ), .B(\ImageBuffer[57][4] ), .C(
        \ImageBuffer[58][4] ), .D(\ImageBuffer[59][4] ), .S0(n4807), .S1(n4811), .Y(n4723) );
  MX4XL U5905 ( .A(\ImageBuffer[40][4] ), .B(\ImageBuffer[41][4] ), .C(
        \ImageBuffer[42][4] ), .D(\ImageBuffer[43][4] ), .S0(n4807), .S1(n4814), .Y(n4728) );
  MX4XL U5906 ( .A(\ImageBuffer[8][4] ), .B(\ImageBuffer[9][4] ), .C(
        \ImageBuffer[10][4] ), .D(\ImageBuffer[11][4] ), .S0(n4802), .S1(n4815), .Y(n4738) );
  MX4XL U5907 ( .A(\ImageBuffer[56][5] ), .B(\ImageBuffer[57][5] ), .C(
        \ImageBuffer[58][5] ), .D(\ImageBuffer[59][5] ), .S0(n4806), .S1(n4815), .Y(n4743) );
  MX4XL U5908 ( .A(\ImageBuffer[40][5] ), .B(\ImageBuffer[41][5] ), .C(
        \ImageBuffer[42][5] ), .D(\ImageBuffer[43][5] ), .S0(N2517), .S1(n4815), .Y(n4748) );
  MX4XL U5909 ( .A(\ImageBuffer[8][5] ), .B(\ImageBuffer[9][5] ), .C(
        \ImageBuffer[10][5] ), .D(\ImageBuffer[11][5] ), .S0(n4804), .S1(n4816), .Y(n4758) );
  MX4XL U5910 ( .A(\ImageBuffer[56][6] ), .B(\ImageBuffer[57][6] ), .C(
        \ImageBuffer[58][6] ), .D(\ImageBuffer[59][6] ), .S0(n4803), .S1(n4816), .Y(n4763) );
  MX4XL U5911 ( .A(\ImageBuffer[40][6] ), .B(\ImageBuffer[41][6] ), .C(
        \ImageBuffer[42][6] ), .D(\ImageBuffer[43][6] ), .S0(n4807), .S1(n4816), .Y(n4768) );
  MX4XL U5912 ( .A(\ImageBuffer[8][6] ), .B(\ImageBuffer[9][6] ), .C(
        \ImageBuffer[10][6] ), .D(\ImageBuffer[11][6] ), .S0(n4808), .S1(n4817), .Y(n4778) );
  MX4XL U5913 ( .A(\ImageBuffer[56][7] ), .B(\ImageBuffer[57][7] ), .C(
        \ImageBuffer[58][7] ), .D(\ImageBuffer[59][7] ), .S0(n4808), .S1(n4817), .Y(n4783) );
  MX4XL U5914 ( .A(\ImageBuffer[40][7] ), .B(\ImageBuffer[41][7] ), .C(
        \ImageBuffer[42][7] ), .D(\ImageBuffer[43][7] ), .S0(n4809), .S1(n4813), .Y(n4788) );
  MX4XL U5915 ( .A(\ImageBuffer[8][7] ), .B(\ImageBuffer[9][7] ), .C(
        \ImageBuffer[10][7] ), .D(\ImageBuffer[11][7] ), .S0(n4809), .S1(n4814), .Y(n4798) );
  MX4XL U5916 ( .A(\ImageBuffer[60][0] ), .B(\ImageBuffer[61][0] ), .C(
        \ImageBuffer[62][0] ), .D(\ImageBuffer[63][0] ), .S0(n4802), .S1(n4811), .Y(n4642) );
  MX4XL U5917 ( .A(\ImageBuffer[44][0] ), .B(\ImageBuffer[45][0] ), .C(
        \ImageBuffer[46][0] ), .D(\ImageBuffer[47][0] ), .S0(n4802), .S1(n4812), .Y(n4647) );
  MX4XL U5918 ( .A(\ImageBuffer[48][0] ), .B(\ImageBuffer[49][0] ), .C(
        \ImageBuffer[50][0] ), .D(\ImageBuffer[51][0] ), .S0(n4802), .S1(n4812), .Y(n4645) );
  MX4XL U5919 ( .A(\ImageBuffer[32][0] ), .B(\ImageBuffer[33][0] ), .C(
        \ImageBuffer[34][0] ), .D(\ImageBuffer[35][0] ), .S0(n4802), .S1(n4814), .Y(n4650) );
  MX4XL U5920 ( .A(\ImageBuffer[52][0] ), .B(\ImageBuffer[53][0] ), .C(
        \ImageBuffer[54][0] ), .D(\ImageBuffer[55][0] ), .S0(n4802), .S1(n4811), .Y(n4644) );
  MX4XL U5921 ( .A(\ImageBuffer[36][0] ), .B(\ImageBuffer[37][0] ), .C(
        \ImageBuffer[38][0] ), .D(\ImageBuffer[39][0] ), .S0(n4802), .S1(n4813), .Y(n4649) );
  MX4XL U5922 ( .A(\ImageBuffer[56][0] ), .B(\ImageBuffer[57][0] ), .C(
        \ImageBuffer[58][0] ), .D(\ImageBuffer[59][0] ), .S0(n4802), .S1(n4811), .Y(n4643) );
  MX4XL U5923 ( .A(\ImageBuffer[40][0] ), .B(\ImageBuffer[41][0] ), .C(
        \ImageBuffer[42][0] ), .D(\ImageBuffer[43][0] ), .S0(n4802), .S1(n4813), .Y(n4648) );
  MX4XL U5924 ( .A(\ImageBuffer[24][0] ), .B(\ImageBuffer[25][0] ), .C(
        \ImageBuffer[26][0] ), .D(\ImageBuffer[27][0] ), .S0(n4802), .S1(n4814), .Y(n4653) );
  MX4XL U5925 ( .A(\ImageBuffer[28][0] ), .B(\ImageBuffer[29][0] ), .C(
        \ImageBuffer[30][0] ), .D(\ImageBuffer[31][0] ), .S0(n4802), .S1(n4814), .Y(n4652) );
  MX4XL U5926 ( .A(\ImageBuffer[20][0] ), .B(\ImageBuffer[21][0] ), .C(
        \ImageBuffer[22][0] ), .D(\ImageBuffer[23][0] ), .S0(n4802), .S1(n4814), .Y(n4654) );
  CLKINVX1 U5927 ( .A(N2517), .Y(n5107) );
  INVX3 U5928 ( .A(n8088), .Y(n8079) );
  CLKBUFX3 U5929 ( .A(N2490), .Y(n3934) );
  CLKBUFX3 U5930 ( .A(n3735), .Y(n3744) );
  INVX6 U5931 ( .A(n7188), .Y(n4860) );
  INVX6 U5932 ( .A(n5046), .Y(n4857) );
  INVX6 U5933 ( .A(n5049), .Y(n4858) );
  AOI222XL U5934 ( .A0(n7306), .A1(n4857), .B0(n7303), .B1(n4860), .C0(n7299), 
        .C1(n4858), .Y(n4851) );
  AOI222XL U5935 ( .A0(n7289), .A1(n4857), .B0(n7288), .B1(n4860), .C0(n7286), 
        .C1(n4858), .Y(n4833) );
  AOI222XL U5936 ( .A0(n7276), .A1(n4857), .B0(n7274), .B1(n4860), .C0(n7271), 
        .C1(n4858), .Y(n4848) );
  AOI222XL U5937 ( .A0(n7262), .A1(n4857), .B0(n7261), .B1(n4860), .C0(n7259), 
        .C1(n4858), .Y(n4832) );
  AOI222XL U5938 ( .A0(n7247), .A1(n4857), .B0(n7246), .B1(n4860), .C0(n7244), 
        .C1(n4858), .Y(n4830) );
  AOI222XL U5939 ( .A0(n7233), .A1(n4857), .B0(n7231), .B1(n4860), .C0(n7228), 
        .C1(n4858), .Y(n4842) );
  AOI222XL U5940 ( .A0(n7217), .A1(n4857), .B0(n7216), .B1(n4860), .C0(n7214), 
        .C1(n4858), .Y(n4828) );
  CLKBUFX3 U5941 ( .A(n3936), .Y(n3940) );
  CLKBUFX3 U5942 ( .A(n5062), .Y(n5056) );
  CLKBUFX3 U5943 ( .A(n5062), .Y(n5055) );
  AOI222XL U5944 ( .A0(n8032), .A1(n4857), .B0(n8026), .B1(n4860), .C0(n8022), 
        .C1(n4858), .Y(n4854) );
  AOI222XL U5945 ( .A0(n8008), .A1(n4857), .B0(n8007), .B1(n4860), .C0(n8005), 
        .C1(n4858), .Y(n4831) );
  AOI222XL U5946 ( .A0(n7985), .A1(n4857), .B0(n7984), .B1(n4860), .C0(n7982), 
        .C1(n4858), .Y(n4829) );
  AOI222XL U5947 ( .A0(n7973), .A1(n4857), .B0(n7972), .B1(n4860), .C0(n7970), 
        .C1(n4858), .Y(n4827) );
  AOI222XL U5948 ( .A0(n7947), .A1(n4857), .B0(n7946), .B1(n4860), .C0(n7944), 
        .C1(n4858), .Y(n4824) );
  AOI222XL U5949 ( .A0(n7933), .A1(n4857), .B0(n7930), .B1(n4860), .C0(n7926), 
        .C1(n4858), .Y(n4856) );
  AOI222XL U5950 ( .A0(n7891), .A1(n4857), .B0(n7889), .B1(n4860), .C0(n7886), 
        .C1(n4858), .Y(n4850) );
  AOI222XL U5951 ( .A0(n7857), .A1(n4857), .B0(n7855), .B1(n4860), .C0(n7852), 
        .C1(n4858), .Y(n4847) );
  AOI222XL U5952 ( .A0(n7831), .A1(n4857), .B0(n7828), .B1(n4860), .C0(n7825), 
        .C1(n4858), .Y(n4841) );
  AOI222XL U5953 ( .A0(n7802), .A1(n4857), .B0(n7801), .B1(n4860), .C0(n7799), 
        .C1(n4858), .Y(n4826) );
  AOI222XL U5954 ( .A0(n7792), .A1(n4857), .B0(n7790), .B1(n4860), .C0(n7787), 
        .C1(n4858), .Y(n4855) );
  AOI222XL U5955 ( .A0(n7768), .A1(n4857), .B0(n7767), .B1(n4860), .C0(n7765), 
        .C1(n4858), .Y(n4823) );
  AOI222XL U5956 ( .A0(n7758), .A1(n4857), .B0(n7756), .B1(n4860), .C0(n7753), 
        .C1(n4858), .Y(n4853) );
  AOI222XL U5957 ( .A0(n7745), .A1(n4857), .B0(n7744), .B1(n4860), .C0(n7742), 
        .C1(n4858), .Y(n4822) );
  AOI222XL U5958 ( .A0(n7732), .A1(n4857), .B0(n7729), .B1(n4860), .C0(n7726), 
        .C1(n4858), .Y(n4852) );
  AOI222XL U5959 ( .A0(n7691), .A1(n4857), .B0(n7689), .B1(n4860), .C0(n7686), 
        .C1(n4858), .Y(n4849) );
  AOI222XL U5960 ( .A0(n7657), .A1(n4857), .B0(n7655), .B1(n4860), .C0(n7652), 
        .C1(n4858), .Y(n4846) );
  AOI222XL U5961 ( .A0(n7631), .A1(n4857), .B0(n7628), .B1(n4860), .C0(n7624), 
        .C1(n4858), .Y(n4840) );
  AOI222XL U5962 ( .A0(n7591), .A1(n4857), .B0(n7589), .B1(n4860), .C0(n7586), 
        .C1(n4858), .Y(n4845) );
  AOI222XL U5963 ( .A0(n7557), .A1(n4857), .B0(n7555), .B1(n4860), .C0(n7552), 
        .C1(n4858), .Y(n4839) );
  AOI222XL U5964 ( .A0(n7531), .A1(n4857), .B0(n7528), .B1(n4860), .C0(n7524), 
        .C1(n4858), .Y(n4836) );
  AOI222XL U5965 ( .A0(n7488), .A1(n4857), .B0(n7486), .B1(n4860), .C0(n7483), 
        .C1(n4858), .Y(n4844) );
  AOI222XL U5966 ( .A0(n7454), .A1(n4857), .B0(n7452), .B1(n4860), .C0(n7449), 
        .C1(n4858), .Y(n4838) );
  AOI222XL U5967 ( .A0(n7428), .A1(n4857), .B0(n7425), .B1(n4860), .C0(n7422), 
        .C1(n4858), .Y(n4835) );
  AOI222XL U5968 ( .A0(n7388), .A1(n4857), .B0(n7386), .B1(n4860), .C0(n7383), 
        .C1(n4858), .Y(n4843) );
  AOI222XL U5969 ( .A0(n7354), .A1(n4857), .B0(n7352), .B1(n4860), .C0(n7349), 
        .C1(n4858), .Y(n4837) );
  AOI222XL U5970 ( .A0(n7328), .A1(n4857), .B0(n7325), .B1(n4860), .C0(n7321), 
        .C1(n4858), .Y(n4834) );
  CLKBUFX3 U5971 ( .A(n5047), .Y(n5048) );
  CLKBUFX3 U5972 ( .A(n7188), .Y(n5047) );
  CLKBUFX3 U5973 ( .A(n6984), .Y(n5031) );
  CLKBUFX3 U5974 ( .A(n6590), .Y(n5005) );
  CLKBUFX3 U5975 ( .A(n6392), .Y(n4992) );
  CLKBUFX3 U5976 ( .A(n6194), .Y(n4980) );
  CLKBUFX3 U5977 ( .A(n5997), .Y(n4967) );
  CLKBUFX3 U5978 ( .A(n6984), .Y(n5032) );
  CLKBUFX3 U5979 ( .A(n6590), .Y(n5006) );
  CLKBUFX3 U5980 ( .A(n5997), .Y(n4968) );
  CLKBUFX3 U5981 ( .A(n5417), .Y(n4954) );
  CLKBUFX3 U5982 ( .A(n4994), .Y(n4993) );
  CLKBUFX3 U5983 ( .A(n5417), .Y(n4955) );
  CLKBUFX3 U5984 ( .A(n5032), .Y(n5033) );
  CLKBUFX3 U5985 ( .A(n6590), .Y(n5007) );
  CLKBUFX3 U5986 ( .A(n6194), .Y(n4981) );
  CLKBUFX3 U5987 ( .A(n5417), .Y(n4956) );
  CLKBUFX3 U5988 ( .A(n6984), .Y(n5034) );
  CLKBUFX3 U5989 ( .A(n5997), .Y(n4969) );
  CLKBUFX3 U5990 ( .A(n4952), .Y(n4951) );
  CLKBUFX3 U5991 ( .A(n5310), .Y(n4952) );
  CLKBUFX3 U5992 ( .A(n4952), .Y(n4953) );
  CLKBUFX3 U5993 ( .A(n6392), .Y(n4994) );
  CLKBUFX3 U5994 ( .A(n6194), .Y(n4982) );
  CLKBUFX3 U5995 ( .A(n7189), .Y(n5049) );
  CLKBUFX3 U5996 ( .A(n5049), .Y(n5050) );
  CLKBUFX3 U5997 ( .A(n5046), .Y(n5045) );
  CLKBUFX3 U5998 ( .A(n5018), .Y(n5019) );
  CLKBUFX3 U5999 ( .A(n5018), .Y(n5020) );
  CLKBUFX3 U6000 ( .A(n5028), .Y(n5029) );
  CLKBUFX3 U6001 ( .A(n6589), .Y(n5002) );
  CLKBUFX3 U6002 ( .A(n4989), .Y(n4990) );
  CLKBUFX3 U6003 ( .A(n4966), .Y(n4963) );
  CLKBUFX3 U6004 ( .A(n5028), .Y(n5030) );
  CLKBUFX3 U6005 ( .A(n4966), .Y(n4964) );
  CLKBUFX3 U6006 ( .A(n6786), .Y(n5015) );
  CLKBUFX3 U6007 ( .A(n4989), .Y(n4991) );
  CLKBUFX3 U6008 ( .A(n6193), .Y(n4977) );
  CLKBUFX3 U6009 ( .A(n6786), .Y(n5016) );
  CLKBUFX3 U6010 ( .A(n6589), .Y(n5004) );
  CLKBUFX3 U6011 ( .A(n6193), .Y(n4978) );
  CLKBUFX3 U6012 ( .A(n4966), .Y(n4965) );
  CLKBUFX3 U6013 ( .A(n6786), .Y(n5017) );
  CLKBUFX3 U6014 ( .A(n6193), .Y(n4979) );
  CLKBUFX3 U6015 ( .A(n3552), .Y(n5021) );
  CLKBUFX3 U6016 ( .A(n6393), .Y(n4995) );
  CLKBUFX3 U6017 ( .A(n6195), .Y(n4983) );
  CLKBUFX3 U6018 ( .A(n4971), .Y(n4970) );
  CLKBUFX3 U6019 ( .A(n5419), .Y(n4957) );
  CLKBUFX3 U6020 ( .A(n5035), .Y(n5036) );
  CLKBUFX3 U6021 ( .A(n5021), .Y(n5022) );
  CLKBUFX3 U6022 ( .A(n5186), .Y(n5008) );
  CLKBUFX3 U6023 ( .A(n6393), .Y(n4996) );
  CLKBUFX3 U6024 ( .A(n6195), .Y(n4984) );
  CLKBUFX3 U6025 ( .A(n5187), .Y(n4971) );
  CLKBUFX3 U6026 ( .A(n5021), .Y(n5023) );
  CLKBUFX3 U6027 ( .A(n5010), .Y(n5009) );
  CLKBUFX3 U6028 ( .A(n6195), .Y(n4985) );
  CLKBUFX3 U6029 ( .A(n4971), .Y(n4972) );
  CLKBUFX3 U6030 ( .A(n5035), .Y(n5037) );
  CLKBUFX3 U6031 ( .A(n6393), .Y(n4997) );
  CLKBUFX3 U6032 ( .A(n5419), .Y(n4958) );
  CLKBUFX3 U6033 ( .A(n5021), .Y(n5024) );
  CLKBUFX3 U6034 ( .A(n5186), .Y(n5010) );
  CLKBUFX3 U6035 ( .A(n4971), .Y(n4973) );
  CLKBUFX3 U6036 ( .A(n5419), .Y(n4959) );
  CLKBUFX3 U6037 ( .A(N2517), .Y(n4803) );
  CLKBUFX3 U6038 ( .A(N2517), .Y(n4804) );
  CLKBUFX3 U6039 ( .A(N2517), .Y(n4805) );
  CLKBUFX3 U6040 ( .A(n5106), .Y(n4806) );
  CLKBUFX3 U6041 ( .A(N2517), .Y(n4807) );
  CLKBUFX3 U6042 ( .A(n5106), .Y(n4808) );
  CLKBUFX3 U6043 ( .A(n4808), .Y(n4809) );
  CLKBUFX3 U6044 ( .A(n4808), .Y(n4802) );
  INVX3 U6045 ( .A(n7609), .Y(n5698) );
  INVX3 U6046 ( .A(n7867), .Y(n5876) );
  INVX3 U6047 ( .A(n7844), .Y(n5858) );
  INVX3 U6048 ( .A(n7810), .Y(n5842) );
  OR2X2 U6049 ( .A(n4908), .B(n7196), .Y(n7526) );
  INVX3 U6050 ( .A(n7866), .Y(n5877) );
  OAI32XL U6051 ( .A0(n7865), .A1(n5053), .A2(n7861), .B0(n5067), .B1(n7829), 
        .Y(n7866) );
  INVX3 U6052 ( .A(n7843), .Y(n5859) );
  INVX3 U6053 ( .A(n7190), .Y(n5418) );
  INVX3 U6054 ( .A(n7195), .Y(n5416) );
  OAI33XL U6055 ( .A0(n7191), .A1(n5053), .A2(n7184), .B0(n7197), .B1(n7194), 
        .B2(n5052), .Y(n7195) );
  INVX3 U6056 ( .A(n7913), .Y(n5913) );
  INVX3 U6057 ( .A(n7900), .Y(n5904) );
  OAI32XL U6058 ( .A0(n7899), .A1(n5053), .A2(n7895), .B0(n5070), .B1(n7829), 
        .Y(n7900) );
  INVX3 U6059 ( .A(n7877), .Y(n5886) );
  OAI32XL U6060 ( .A0(n7876), .A1(n5053), .A2(n7872), .B0(n5068), .B1(n7829), 
        .Y(n7877) );
  INVX3 U6061 ( .A(n7814), .Y(n5841) );
  INVX3 U6062 ( .A(n7778), .Y(n5814) );
  INVX3 U6063 ( .A(n7714), .Y(n5769) );
  INVX3 U6064 ( .A(n7700), .Y(n5760) );
  OAI32XL U6065 ( .A0(n7699), .A1(n5053), .A2(n7695), .B0(n5070), .B1(n7629), 
        .Y(n7700) );
  INVX3 U6066 ( .A(n7677), .Y(n5742) );
  OAI32XL U6067 ( .A0(n7676), .A1(n5053), .A2(n7672), .B0(n5068), .B1(n7629), 
        .Y(n7677) );
  INVX3 U6068 ( .A(n7666), .Y(n5733) );
  INVX3 U6069 ( .A(n7643), .Y(n5715) );
  INVX3 U6070 ( .A(n7613), .Y(n5697) );
  OAI33XL U6071 ( .A0(n7610), .A1(n5053), .A2(n7606), .B0(n7529), .B1(n7611), 
        .B2(n5071), .Y(n7613) );
  INVX3 U6072 ( .A(n7600), .Y(n5688) );
  OAI32XL U6073 ( .A0(n7599), .A1(n5053), .A2(n7595), .B0(n5070), .B1(n7529), 
        .Y(n7600) );
  INVX3 U6074 ( .A(n7577), .Y(n5670) );
  OAI32XL U6075 ( .A0(n7576), .A1(n5053), .A2(n7572), .B0(n5068), .B1(n7529), 
        .Y(n7577) );
  INVX3 U6076 ( .A(n7566), .Y(n5661) );
  OAI32XL U6077 ( .A0(n7565), .A1(n5053), .A2(n7561), .B0(n5067), .B1(n7529), 
        .Y(n7566) );
  INVX3 U6078 ( .A(n7543), .Y(n5643) );
  OAI32XL U6079 ( .A0(n7542), .A1(n5053), .A2(n7538), .B0(n8057), .B1(n7529), 
        .Y(n7543) );
  INVX3 U6080 ( .A(n7512), .Y(n5625) );
  INVX3 U6081 ( .A(n7497), .Y(n5616) );
  OAI32XL U6082 ( .A0(n7496), .A1(n5053), .A2(n7492), .B0(n5070), .B1(n7426), 
        .Y(n7497) );
  INVX3 U6083 ( .A(n7474), .Y(n5598) );
  OAI32XL U6084 ( .A0(n7473), .A1(n5053), .A2(n7469), .B0(n5068), .B1(n7426), 
        .Y(n7474) );
  INVX3 U6085 ( .A(n7463), .Y(n5589) );
  OAI32XL U6086 ( .A0(n7462), .A1(n5053), .A2(n7458), .B0(n5067), .B1(n7426), 
        .Y(n7463) );
  INVX3 U6087 ( .A(n7440), .Y(n5571) );
  OAI32XL U6088 ( .A0(n7439), .A1(n5053), .A2(n7435), .B0(n8057), .B1(n7426), 
        .Y(n7440) );
  INVX3 U6089 ( .A(n7411), .Y(n5553) );
  INVX3 U6090 ( .A(n7397), .Y(n5544) );
  INVX3 U6091 ( .A(n7374), .Y(n5526) );
  INVX3 U6092 ( .A(n7363), .Y(n5517) );
  INVX3 U6093 ( .A(n7340), .Y(n5499) );
  CLKBUFX3 U6094 ( .A(n5063), .Y(n5054) );
  CLKBUFX3 U6095 ( .A(n5064), .Y(n5063) );
  CLKBUFX3 U6096 ( .A(n5118), .Y(n4121) );
  CLKBUFX3 U6097 ( .A(n5118), .Y(n3746) );
  CLKBUFX3 U6098 ( .A(n5118), .Y(n4120) );
  INVX3 U6099 ( .A(n7864), .Y(n5878) );
  OAI32XL U6100 ( .A0(n7865), .A1(n7192), .A2(n7861), .B0(n5067), .B1(n3369), 
        .Y(n7864) );
  INVX3 U6101 ( .A(n7841), .Y(n5860) );
  OAI32XL U6102 ( .A0(n7842), .A1(n7192), .A2(n7838), .B0(n8057), .B1(n3369), 
        .Y(n7841) );
  CLKBUFX3 U6103 ( .A(N2495), .Y(n3759) );
  CLKBUFX3 U6104 ( .A(N2513), .Y(n4640) );
  CLKBUFX3 U6105 ( .A(n4135), .Y(n4136) );
  INVX3 U6106 ( .A(n5103), .Y(n5101) );
  CLKBUFX6 U6107 ( .A(n3944), .Y(n5081) );
  INVX6 U6108 ( .A(n5087), .Y(n5083) );
  CLKBUFX3 U6109 ( .A(n3549), .Y(n5067) );
  INVX6 U6110 ( .A(n5097), .Y(n5094) );
  INVX6 U6111 ( .A(n5102), .Y(n5099) );
  CLKBUFX3 U6112 ( .A(n3547), .Y(n5065) );
  CLKBUFX3 U6113 ( .A(n5044), .Y(n5043) );
  CLKBUFX3 U6114 ( .A(n5248), .Y(n4966) );
  INVX3 U6115 ( .A(n8057), .Y(n7210) );
  CLKBUFX6 U6116 ( .A(n3944), .Y(n5082) );
  CLKBUFX6 U6117 ( .A(n5074), .Y(n5073) );
  INVX6 U6118 ( .A(n5086), .Y(n5084) );
  INVX6 U6119 ( .A(n5097), .Y(n5095) );
  INVX6 U6120 ( .A(n5102), .Y(n5100) );
  CLKBUFX3 U6121 ( .A(n5043), .Y(n5042) );
  CLKBUFX3 U6122 ( .A(n3548), .Y(n5052) );
  CLKBUFX3 U6123 ( .A(N2518), .Y(n4811) );
  CLKBUFX3 U6124 ( .A(N2518), .Y(n4812) );
  CLKBUFX3 U6125 ( .A(N2518), .Y(n4813) );
  CLKBUFX3 U6126 ( .A(N2518), .Y(n4814) );
  CLKBUFX3 U6127 ( .A(n4810), .Y(n4815) );
  CLKBUFX3 U6128 ( .A(n4810), .Y(n4816) );
  CLKBUFX3 U6129 ( .A(n4810), .Y(n4817) );
  OAI2BB2X2 U6130 ( .B0(n7180), .B1(n3344), .A0N(n5401), .A1N(N2538), .Y(n5411) );
  CLKXOR2X4 U6131 ( .A(n5125), .B(n5127), .Y(N2497) );
  CLKXOR2X4 U6132 ( .A(n5125), .B(\add_80/carry[4] ), .Y(N2503) );
  AOI211X1 U6133 ( .A0(n5150), .A1(n5149), .B0(n5148), .C0(n5147), .Y(n5152)
         );
  CLKBUFX3 U6134 ( .A(n5080), .Y(n5078) );
  CLKBUFX3 U6135 ( .A(n5982), .Y(n4945) );
  CLKBUFX3 U6136 ( .A(n5981), .Y(n4942) );
  CLKBUFX3 U6137 ( .A(n5945), .Y(n4938) );
  CLKBUFX3 U6138 ( .A(n5127), .Y(n3733) );
  CLKBUFX3 U6139 ( .A(n5954), .Y(n4939) );
  CLKBUFX3 U6140 ( .A(n5918), .Y(n4935) );
  OAI22XL U6141 ( .A0(n7315), .A1(n7918), .B0(n7919), .B1(n3344), .Y(n5918) );
  CLKINVX1 U6142 ( .A(n4868), .Y(n5278) );
  CLKINVX1 U6143 ( .A(n4868), .Y(n5248) );
  CLKINVX1 U6144 ( .A(n4873), .Y(n5308) );
  CLKINVX1 U6145 ( .A(n4873), .Y(n5276) );
  CLKINVX1 U6146 ( .A(n4873), .Y(n5247) );
  CLKBUFX3 U6147 ( .A(n3366), .Y(n5064) );
  AOI222XL U6148 ( .A0(n7961), .A1(N2765), .B0(n7959), .B1(n4860), .C0(n7956), 
        .C1(N2781), .Y(n4859) );
  CLKINVX1 U6149 ( .A(n4867), .Y(n5250) );
  CLKINVX1 U6150 ( .A(n4867), .Y(n5310) );
  CLKINVX1 U6151 ( .A(n4862), .Y(n5219) );
  CLKINVX1 U6152 ( .A(n4862), .Y(n5187) );
  CLKINVX1 U6153 ( .A(n4861), .Y(n5157) );
  CLKINVX1 U6154 ( .A(n4861), .Y(n5188) );
  CLKBUFX3 U6155 ( .A(N2513), .Y(n4641) );
  CLKBUFX3 U6156 ( .A(n7734), .Y(n4926) );
  NAND3X2 U6157 ( .A(n7515), .B(n7717), .C(n5127), .Y(n7935) );
  CLKBUFX3 U6158 ( .A(n7533), .Y(n4908) );
  NAND3XL U6159 ( .A(N2498), .B(n7515), .C(n5127), .Y(n7533) );
  CLKBUFX3 U6160 ( .A(n6586), .Y(n4998) );
  CLKBUFX3 U6161 ( .A(n6388), .Y(n4986) );
  CLKBUFX3 U6162 ( .A(n6980), .Y(n5025) );
  CLKBUFX3 U6163 ( .A(n6783), .Y(n5011) );
  CLKBUFX3 U6164 ( .A(n6388), .Y(n4987) );
  CLKBUFX3 U6165 ( .A(n5410), .Y(n4948) );
  CLKBUFX3 U6166 ( .A(n6783), .Y(n5012) );
  CLKBUFX3 U6167 ( .A(n6586), .Y(n4999) );
  CLKBUFX3 U6168 ( .A(n6190), .Y(n4974) );
  CLKBUFX3 U6169 ( .A(n5994), .Y(n4960) );
  CLKBUFX3 U6170 ( .A(n5410), .Y(n4949) );
  CLKBUFX3 U6171 ( .A(n7178), .Y(n5038) );
  CLKBUFX3 U6172 ( .A(n6980), .Y(n5026) );
  CLKBUFX3 U6173 ( .A(n6783), .Y(n5013) );
  CLKBUFX3 U6174 ( .A(n6586), .Y(n5000) );
  CLKBUFX3 U6175 ( .A(n6388), .Y(n4988) );
  CLKBUFX3 U6176 ( .A(n6190), .Y(n4975) );
  CLKBUFX3 U6177 ( .A(n5994), .Y(n4961) );
  CLKBUFX3 U6178 ( .A(n5410), .Y(n4950) );
  CLKBUFX3 U6179 ( .A(n7178), .Y(n5039) );
  CLKBUFX3 U6180 ( .A(n6980), .Y(n5027) );
  CLKBUFX3 U6181 ( .A(n6783), .Y(n5014) );
  CLKBUFX3 U6182 ( .A(n6586), .Y(n5001) );
  CLKBUFX3 U6183 ( .A(n6190), .Y(n4976) );
  CLKBUFX3 U6184 ( .A(n5994), .Y(n4962) );
  CLKBUFX3 U6185 ( .A(n3946), .Y(n5089) );
  CLKBUFX3 U6186 ( .A(n7178), .Y(n5040) );
  CLKBUFX3 U6187 ( .A(n3559), .Y(n5070) );
  CLKBUFX3 U6188 ( .A(n3560), .Y(n5068) );
  CLKBUFX3 U6189 ( .A(n3562), .Y(n5069) );
  CLKBUFX3 U6190 ( .A(n3561), .Y(n5066) );
  CLKBUFX3 U6191 ( .A(n7330), .Y(n4890) );
  CLKBUFX3 U6192 ( .A(n6787), .Y(n5018) );
  CLKBUFX3 U6193 ( .A(n6983), .Y(n5028) );
  CLKBUFX3 U6194 ( .A(n6985), .Y(n5035) );
  CLKBUFX3 U6195 ( .A(n6391), .Y(n4989) );
  CLKBUFX3 U6196 ( .A(n5041), .Y(n5044) );
  CLKBUFX3 U6197 ( .A(n3558), .Y(n5071) );
  CLKBUFX3 U6198 ( .A(n5105), .Y(n4810) );
  CLKBUFX3 U6199 ( .A(N2520), .Y(n4820) );
  CLKBUFX3 U6200 ( .A(n5104), .Y(n4821) );
  CLKBUFX3 U6201 ( .A(N2519), .Y(n4818) );
  CLKBUFX3 U6202 ( .A(N2519), .Y(n4819) );
  MX4X1 U6203 ( .A(n4265), .B(n4263), .C(n4264), .D(n4262), .S0(n5108), .S1(
        n3487), .Y(n4266) );
  MX4X1 U6204 ( .A(n4275), .B(n4273), .C(n4274), .D(n4272), .S0(n5108), .S1(
        n3487), .Y(n4276) );
  MX4X1 U6205 ( .A(n4260), .B(n4258), .C(n4259), .D(n4257), .S0(n5108), .S1(
        n3487), .Y(n4261) );
  MX4X1 U6206 ( .A(n4160), .B(n4158), .C(n4159), .D(n4157), .S0(n5108), .S1(
        n3487), .Y(n4161) );
  MX4X1 U6207 ( .A(n4165), .B(n4163), .C(n4164), .D(n4162), .S0(n5108), .S1(
        n3487), .Y(n4166) );
  MX4X1 U6208 ( .A(n4170), .B(n4168), .C(n4169), .D(n4167), .S0(n5108), .S1(
        n3487), .Y(n4171) );
  OAI22XL U6209 ( .A0(n7293), .A1(n7720), .B0(n7806), .B1(n3344), .Y(n5837) );
  MX4X1 U6210 ( .A(n3581), .B(n3579), .C(n3580), .D(n3578), .S0(n3733), .S1(
        n3758), .Y(n3582) );
  MX4X1 U6211 ( .A(n3576), .B(n3574), .C(n3575), .D(n3573), .S0(n3733), .S1(
        n3758), .Y(n3577) );
  MX4X1 U6212 ( .A(n4517), .B(n4515), .C(n4516), .D(n4514), .S0(n3496), .S1(
        n4639), .Y(n4518) );
  MX4X1 U6213 ( .A(n4507), .B(n4505), .C(n4506), .D(n4504), .S0(n3496), .S1(
        n4641), .Y(n4508) );
  MX4X1 U6214 ( .A(n4512), .B(n4510), .C(n4511), .D(n4509), .S0(n3496), .S1(
        n4639), .Y(n4513) );
  MX4X1 U6215 ( .A(n4417), .B(n4415), .C(n4416), .D(n4414), .S0(n3503), .S1(
        n3495), .Y(n4418) );
  MX4X1 U6216 ( .A(n4427), .B(n4425), .C(n4426), .D(n4424), .S0(n3503), .S1(
        n3495), .Y(n4428) );
  MX4X1 U6217 ( .A(n4422), .B(n4420), .C(n4421), .D(n4419), .S0(n3503), .S1(
        n3495), .Y(n4423) );
  MXI4X4 U6218 ( .A(n3779), .B(n3769), .C(n3774), .D(n3764), .S0(N2492), .S1(
        N2491), .Y(n3572) );
  MX4X1 U6219 ( .A(n3612), .B(n3602), .C(n3607), .D(n3597), .S0(n4946), .S1(
        n5125), .Y(N2780) );
  MX4X1 U6220 ( .A(n3601), .B(n3599), .C(n3600), .D(n3598), .S0(n3733), .S1(
        n3759), .Y(n3602) );
  MX4X1 U6221 ( .A(n3631), .B(n3629), .C(n3630), .D(n3628), .S0(n3734), .S1(
        n3758), .Y(n3632) );
  MX4X1 U6222 ( .A(n3621), .B(n3619), .C(n3620), .D(n3618), .S0(n3734), .S1(
        n3758), .Y(n3622) );
  MX4X1 U6223 ( .A(n3672), .B(n3662), .C(n3667), .D(n3657), .S0(n4946), .S1(
        n5125), .Y(N2777) );
  MX4X1 U6224 ( .A(n3671), .B(n3669), .C(n3670), .D(n3668), .S0(n3734), .S1(
        n3759), .Y(n3672) );
  MX4X1 U6225 ( .A(n3661), .B(n3659), .C(n3660), .D(n3658), .S0(n3734), .S1(
        n3758), .Y(n3662) );
  MX4X1 U6226 ( .A(n3652), .B(n3642), .C(n3647), .D(n3637), .S0(n4946), .S1(
        n5125), .Y(N2778) );
  MX4X1 U6227 ( .A(n3651), .B(n3649), .C(n3650), .D(n3648), .S0(n3734), .S1(
        n3758), .Y(n3652) );
  MX4X1 U6228 ( .A(n3828), .B(n3826), .C(n3827), .D(n3825), .S0(n3933), .S1(
        n3409), .Y(n3829) );
  CLKBUFX3 U6229 ( .A(n5972), .Y(n4941) );
  OAI22XL U6230 ( .A0(n7280), .A1(n7918), .B0(n8001), .B1(n3344), .Y(n5972) );
  CLKBUFX3 U6231 ( .A(n5936), .Y(n4937) );
  OAI22XL U6232 ( .A0(n7222), .A1(n7918), .B0(n7951), .B1(n3344), .Y(n5936) );
  CLKBUFX3 U6233 ( .A(n5909), .Y(n4934) );
  CLKBUFX3 U6234 ( .A(n5900), .Y(n4933) );
  OAI22XL U6235 ( .A0(n7280), .A1(n7819), .B0(n7894), .B1(n3344), .Y(n5900) );
  CLKBUFX3 U6236 ( .A(n5873), .Y(n4930) );
  CLKBUFX3 U6237 ( .A(n5864), .Y(n4929) );
  OAI22XL U6238 ( .A0(n7222), .A1(n7819), .B0(n7848), .B1(n3344), .Y(n5864) );
  CLKBUFX3 U6239 ( .A(n5828), .Y(n4924) );
  OAI22XL U6240 ( .A0(n7280), .A1(n7720), .B0(n7795), .B1(n3344), .Y(n5828) );
  CLKBUFX3 U6241 ( .A(n5801), .Y(n4921) );
  CLKBUFX3 U6242 ( .A(n5792), .Y(n4920) );
  OAI22XL U6243 ( .A0(n7222), .A1(n7720), .B0(n7749), .B1(n3344), .Y(n5792) );
  CLKBUFX3 U6244 ( .A(n5765), .Y(n4916) );
  OAI22XL U6245 ( .A0(n7293), .A1(n7618), .B0(n7705), .B1(n3344), .Y(n5765) );
  CLKBUFX3 U6246 ( .A(n5756), .Y(n4915) );
  OAI22XL U6247 ( .A0(n7280), .A1(n7618), .B0(n7694), .B1(n3344), .Y(n5756) );
  CLKBUFX3 U6248 ( .A(n5729), .Y(n4912) );
  OAI22XL U6249 ( .A0(n7238), .A1(n7618), .B0(n7660), .B1(n3344), .Y(n5729) );
  CLKBUFX3 U6250 ( .A(n5720), .Y(n4911) );
  OAI22XL U6251 ( .A0(n7222), .A1(n7618), .B0(n7648), .B1(n3344), .Y(n5720) );
  CLKBUFX3 U6252 ( .A(n5693), .Y(n4907) );
  CLKBUFX3 U6253 ( .A(n5684), .Y(n4906) );
  OAI22XL U6254 ( .A0(n7280), .A1(n7518), .B0(n7594), .B1(n3344), .Y(n5684) );
  CLKBUFX3 U6255 ( .A(n5657), .Y(n4903) );
  CLKBUFX3 U6256 ( .A(n5648), .Y(n4902) );
  OAI22XL U6257 ( .A0(n7222), .A1(n7518), .B0(n7548), .B1(n3344), .Y(n5648) );
  CLKBUFX3 U6258 ( .A(n5621), .Y(n4898) );
  CLKBUFX3 U6259 ( .A(n5612), .Y(n4897) );
  OAI22XL U6260 ( .A0(n7280), .A1(n7416), .B0(n7491), .B1(n3344), .Y(n5612) );
  CLKBUFX3 U6261 ( .A(n5585), .Y(n4894) );
  CLKBUFX3 U6262 ( .A(n5576), .Y(n4893) );
  OAI22XL U6263 ( .A0(n7222), .A1(n7416), .B0(n7445), .B1(n3344), .Y(n5576) );
  CLKBUFX3 U6264 ( .A(n5549), .Y(n4889) );
  CLKBUFX3 U6265 ( .A(n5540), .Y(n4888) );
  OAI22XL U6266 ( .A0(n7280), .A1(n7314), .B0(n7391), .B1(n3344), .Y(n5540) );
  CLKBUFX3 U6267 ( .A(n5513), .Y(n4885) );
  OAI22XL U6268 ( .A0(n7238), .A1(n7314), .B0(n7357), .B1(n3344), .Y(n5513) );
  CLKBUFX3 U6269 ( .A(n5504), .Y(n4884) );
  OAI22XL U6270 ( .A0(n7222), .A1(n7314), .B0(n7345), .B1(n3344), .Y(n5504) );
  CLKBUFX3 U6271 ( .A(n5963), .Y(n4940) );
  OAI22XL U6272 ( .A0(n7266), .A1(n7918), .B0(n7989), .B1(n3344), .Y(n5963) );
  CLKBUFX3 U6273 ( .A(n5927), .Y(n4936) );
  OAI22XL U6274 ( .A0(n7208), .A1(n7918), .B0(n7939), .B1(n3344), .Y(n5927) );
  CLKBUFX3 U6275 ( .A(n5891), .Y(n4932) );
  OAI22XL U6276 ( .A0(n7266), .A1(n7819), .B0(n7882), .B1(n3344), .Y(n5891) );
  CLKBUFX3 U6277 ( .A(n5855), .Y(n4928) );
  OAI22XL U6278 ( .A0(n7208), .A1(n7819), .B0(n7837), .B1(n3344), .Y(n5855) );
  CLKBUFX3 U6279 ( .A(n5819), .Y(n4923) );
  OAI22XL U6280 ( .A0(n7266), .A1(n7720), .B0(n7783), .B1(n3344), .Y(n5819) );
  CLKBUFX3 U6281 ( .A(n5783), .Y(n4919) );
  OAI22XL U6282 ( .A0(n7208), .A1(n7720), .B0(n7738), .B1(n3344), .Y(n5783) );
  CLKBUFX3 U6283 ( .A(n5747), .Y(n4914) );
  OAI22XL U6284 ( .A0(n7266), .A1(n7618), .B0(n7682), .B1(n3344), .Y(n5747) );
  CLKBUFX3 U6285 ( .A(n5711), .Y(n4910) );
  OAI22XL U6286 ( .A0(n7208), .A1(n7618), .B0(n7637), .B1(n3344), .Y(n5711) );
  CLKBUFX3 U6287 ( .A(n5675), .Y(n4905) );
  OAI22XL U6288 ( .A0(n7266), .A1(n7518), .B0(n7582), .B1(n3344), .Y(n5675) );
  CLKBUFX3 U6289 ( .A(n5639), .Y(n4901) );
  OAI22XL U6290 ( .A0(n7208), .A1(n7518), .B0(n7537), .B1(n3344), .Y(n5639) );
  CLKBUFX3 U6291 ( .A(n5603), .Y(n4896) );
  OAI22XL U6292 ( .A0(n7266), .A1(n7416), .B0(n7479), .B1(n3344), .Y(n5603) );
  CLKBUFX3 U6293 ( .A(n5567), .Y(n4892) );
  OAI22XL U6294 ( .A0(n7208), .A1(n7416), .B0(n7434), .B1(n3344), .Y(n5567) );
  CLKBUFX3 U6295 ( .A(n5531), .Y(n4887) );
  OAI22XL U6296 ( .A0(n7266), .A1(n7314), .B0(n7379), .B1(n3344), .Y(n5531) );
  CLKBUFX3 U6297 ( .A(n5495), .Y(n4883) );
  OAI22XL U6298 ( .A0(n7208), .A1(n7314), .B0(n7334), .B1(n3344), .Y(n5495) );
  CLKBUFX3 U6299 ( .A(n5486), .Y(n4882) );
  OAI22XL U6300 ( .A0(n7314), .A1(n7315), .B0(n7316), .B1(n3344), .Y(n5486) );
  CLKBUFX3 U6301 ( .A(n5128), .Y(n4110) );
  CLKBUFX3 U6302 ( .A(n5477), .Y(n4880) );
  OAI22XL U6303 ( .A0(n7207), .A1(n7293), .B0(n7294), .B1(n3344), .Y(n5477) );
  CLKBUFX3 U6304 ( .A(n5468), .Y(n4879) );
  OAI22XL U6305 ( .A0(n7207), .A1(n7280), .B0(n7281), .B1(n3344), .Y(n5468) );
  CLKBUFX3 U6306 ( .A(n5459), .Y(n4878) );
  OAI22XL U6307 ( .A0(n7207), .A1(n7266), .B0(n7267), .B1(n3344), .Y(n5459) );
  CLKBUFX3 U6308 ( .A(n5450), .Y(n4877) );
  OAI22XL U6309 ( .A0(n7207), .A1(n7253), .B0(n7254), .B1(n3344), .Y(n5450) );
  CLKBUFX3 U6310 ( .A(n5441), .Y(n4876) );
  OAI22XL U6311 ( .A0(n7207), .A1(n7238), .B0(n7239), .B1(n3344), .Y(n5441) );
  CLKBUFX3 U6312 ( .A(n5432), .Y(n4875) );
  OAI22XL U6313 ( .A0(n7207), .A1(n7222), .B0(n7223), .B1(n3344), .Y(n5432) );
  CLKBUFX3 U6314 ( .A(n5423), .Y(n4874) );
  OAI22XL U6315 ( .A0(n7207), .A1(n7208), .B0(n7209), .B1(n3344), .Y(n5423) );
  CLKBUFX3 U6316 ( .A(n5882), .Y(n4931) );
  CLKBUFX3 U6317 ( .A(n5810), .Y(n4922) );
  CLKBUFX3 U6318 ( .A(n5738), .Y(n4913) );
  OAI22XL U6319 ( .A0(n7253), .A1(n7618), .B0(n7671), .B1(n3344), .Y(n5738) );
  CLKBUFX3 U6320 ( .A(n5666), .Y(n4904) );
  OAI22XL U6321 ( .A0(n7253), .A1(n7518), .B0(n7571), .B1(n3344), .Y(n5666) );
  CLKBUFX3 U6322 ( .A(n5594), .Y(n4895) );
  CLKBUFX3 U6323 ( .A(n5522), .Y(n4886) );
  OAI22XL U6324 ( .A0(n7253), .A1(n7314), .B0(n7368), .B1(n3344), .Y(n5522) );
  CLKBUFX3 U6325 ( .A(n5846), .Y(n4927) );
  OAI22XL U6326 ( .A0(n7315), .A1(n7819), .B0(n7820), .B1(n3344), .Y(n5846) );
  CLKBUFX3 U6327 ( .A(n5774), .Y(n4918) );
  OAI22XL U6328 ( .A0(n7315), .A1(n7720), .B0(n7721), .B1(n3344), .Y(n5774) );
  CLKBUFX3 U6329 ( .A(n5702), .Y(n4909) );
  OAI22XL U6330 ( .A0(n7315), .A1(n7618), .B0(n7619), .B1(n3344), .Y(n5702) );
  CLKBUFX3 U6331 ( .A(n5630), .Y(n4900) );
  OAI22XL U6332 ( .A0(n7315), .A1(n7518), .B0(n7519), .B1(n3344), .Y(n5630) );
  CLKBUFX3 U6333 ( .A(n5558), .Y(n4891) );
  OAI22XL U6334 ( .A0(n7315), .A1(n7416), .B0(n7417), .B1(n3344), .Y(n5558) );
  AND2X2 U6335 ( .A(n5127), .B(n5125), .Y(\add_79/carry[5] ) );
  MX4X1 U6336 ( .A(n4036), .B(n4034), .C(n4035), .D(n4033), .S0(n4108), .S1(
        n4135), .Y(n4037) );
  CLKINVX1 U6337 ( .A(n3948), .Y(n5098) );
  MX4X1 U6338 ( .A(n4087), .B(n4077), .C(n4082), .D(n4072), .S0(N2498), .S1(
        N2497), .Y(n3948) );
  MX4X1 U6339 ( .A(n4086), .B(n4084), .C(n4085), .D(n4083), .S0(n4109), .S1(
        n4136), .Y(n4087) );
  MX4X1 U6340 ( .A(n4027), .B(n4017), .C(n4022), .D(n4012), .S0(N2498), .S1(
        N2497), .Y(n3945) );
  MX4X1 U6341 ( .A(n4026), .B(n4024), .C(n4025), .D(n4023), .S0(n4108), .S1(
        n4135), .Y(n4027) );
  MX4X1 U6342 ( .A(n3692), .B(n3682), .C(n3687), .D(n3677), .S0(n4946), .S1(
        n5125), .Y(N2776) );
  MX4X1 U6343 ( .A(n3691), .B(n3689), .C(n3690), .D(n3688), .S0(n3734), .S1(
        n3759), .Y(n3692) );
  MX4X1 U6344 ( .A(n3681), .B(n3679), .C(n3680), .D(n3678), .S0(n3734), .S1(
        n3759), .Y(n3682) );
  MX4X1 U6345 ( .A(n3732), .B(n3722), .C(n3727), .D(n3717), .S0(n4946), .S1(
        n5125), .Y(N2774) );
  CLKINVX1 U6346 ( .A(n3949), .Y(n5103) );
  MX4X1 U6347 ( .A(n4107), .B(n4097), .C(n4102), .D(n4092), .S0(N2498), .S1(
        N2497), .Y(n3949) );
  MX4X1 U6348 ( .A(n4106), .B(n4104), .C(n4105), .D(n4103), .S0(n4109), .S1(
        n4136), .Y(n4107) );
  CLKBUFX3 U6349 ( .A(n7430), .Y(n4899) );
  NAND3XL U6350 ( .A(n5128), .B(n7515), .C(N2498), .Y(n7430) );
  CLKBUFX3 U6351 ( .A(n7633), .Y(n4917) );
  NAND3XL U6352 ( .A(n5128), .B(n7717), .C(N2497), .Y(n7633) );
  CLKBUFX3 U6353 ( .A(n7202), .Y(n4881) );
  BUFX16 U6354 ( .A(N2541), .Y(IRAM_valid) );
  CLKBUFX3 U6355 ( .A(n7179), .Y(n5041) );
  ADDHXL U6356 ( .A(N2519), .B(\add_134/carry[2] ), .CO(\add_134/carry[3] ), 
        .S(N2569) );
  ADDHXL U6357 ( .A(n5104), .B(\add_134/carry[3] ), .CO(\add_134/carry[4] ), 
        .S(N2570) );
  ADDHXL U6358 ( .A(n5105), .B(n5106), .CO(\add_134/carry[2] ), .S(N2568) );
  CLKINVX1 U6359 ( .A(n4859), .Y(n7955) );
  CLKINVX1 U6360 ( .A(n4856), .Y(n7925) );
  CLKINVX1 U6361 ( .A(n4850), .Y(n7885) );
  CLKINVX1 U6362 ( .A(n4847), .Y(n7851) );
  CLKINVX1 U6363 ( .A(n4841), .Y(n7824) );
  CLKINVX1 U6364 ( .A(n4855), .Y(n7786) );
  CLKINVX1 U6365 ( .A(n4853), .Y(n7752) );
  CLKINVX1 U6366 ( .A(n4852), .Y(n7725) );
  CLKINVX1 U6367 ( .A(n4849), .Y(n7685) );
  CLKINVX1 U6368 ( .A(n4846), .Y(n7651) );
  CLKINVX1 U6369 ( .A(n4840), .Y(n7623) );
  CLKINVX1 U6370 ( .A(n4845), .Y(n7585) );
  CLKINVX1 U6371 ( .A(n4839), .Y(n7551) );
  CLKINVX1 U6372 ( .A(n4836), .Y(n7523) );
  CLKINVX1 U6373 ( .A(n4844), .Y(n7482) );
  CLKINVX1 U6374 ( .A(n4838), .Y(n7448) );
  CLKINVX1 U6375 ( .A(n4835), .Y(n7421) );
  CLKINVX1 U6376 ( .A(n4843), .Y(n7382) );
  CLKINVX1 U6377 ( .A(n4837), .Y(n7348) );
  CLKINVX1 U6378 ( .A(n4834), .Y(n7320) );
  CLKINVX1 U6379 ( .A(n4851), .Y(n7298) );
  CLKINVX1 U6380 ( .A(n4848), .Y(n7270) );
  CLKINVX1 U6381 ( .A(n4842), .Y(n7227) );
  CLKINVX1 U6382 ( .A(n4854), .Y(n8019) );
  CLKINVX1 U6383 ( .A(n4831), .Y(n8004) );
  CLKINVX1 U6384 ( .A(n4829), .Y(n7981) );
  CLKINVX1 U6385 ( .A(n4827), .Y(n7969) );
  CLKINVX1 U6386 ( .A(n4824), .Y(n7943) );
  OAI222XL U6387 ( .A0(n5858), .A1(n5045), .B0(n5859), .B1(n5047), .C0(n5860), 
        .C1(n5050), .Y(n7840) );
  CLKINVX1 U6388 ( .A(n4826), .Y(n7798) );
  CLKINVX1 U6389 ( .A(n4823), .Y(n7764) );
  CLKINVX1 U6390 ( .A(n4822), .Y(n7741) );
  CLKINVX1 U6391 ( .A(n4833), .Y(n7285) );
  CLKINVX1 U6392 ( .A(n4832), .Y(n7258) );
  CLKINVX1 U6393 ( .A(n4830), .Y(n7243) );
  CLKINVX1 U6394 ( .A(n4828), .Y(n7213) );
  MX4X1 U6395 ( .A(\ImageBuffer[16][3] ), .B(\ImageBuffer[17][3] ), .C(
        \ImageBuffer[18][3] ), .D(\ImageBuffer[19][3] ), .S0(n3935), .S1(n4312), .Y(n4210) );
  MX4X1 U6396 ( .A(\ImageBuffer[24][3] ), .B(\ImageBuffer[25][3] ), .C(
        \ImageBuffer[26][3] ), .D(\ImageBuffer[27][3] ), .S0(n3935), .S1(n4309), .Y(n4208) );
  MX4X1 U6397 ( .A(\ImageBuffer[20][3] ), .B(\ImageBuffer[21][3] ), .C(
        \ImageBuffer[22][3] ), .D(\ImageBuffer[23][3] ), .S0(n4298), .S1(n4305), .Y(n4209) );
  OAI21XL U6398 ( .A0(n6917), .A1(n5808), .B0(n6918), .Y(n8454) );
  OAI21XL U6399 ( .A0(n6899), .A1(n5754), .B0(n6900), .Y(n8448) );
  OAI21XL U6400 ( .A0(n6926), .A1(n5835), .B0(n6927), .Y(n8457) );
  MX4X1 U6401 ( .A(\ImageBuffer[20][3] ), .B(\ImageBuffer[21][3] ), .C(
        \ImageBuffer[22][3] ), .D(\ImageBuffer[23][3] ), .S0(n3513), .S1(n3473), .Y(n4391) );
  MX4X1 U6402 ( .A(\ImageBuffer[52][3] ), .B(\ImageBuffer[53][3] ), .C(
        \ImageBuffer[54][3] ), .D(\ImageBuffer[55][3] ), .S0(n3521), .S1(n3473), .Y(n4381) );
  MX4X1 U6403 ( .A(\ImageBuffer[36][2] ), .B(\ImageBuffer[37][2] ), .C(
        \ImageBuffer[38][2] ), .D(\ImageBuffer[39][2] ), .S0(n3740), .S1(n4124), .Y(n3995) );
  MX4X1 U6404 ( .A(\ImageBuffer[4][2] ), .B(\ImageBuffer[5][2] ), .C(
        \ImageBuffer[6][2] ), .D(\ImageBuffer[7][2] ), .S0(n3740), .S1(n3754), 
        .Y(n4005) );
  MX4X1 U6405 ( .A(\ImageBuffer[36][0] ), .B(\ImageBuffer[37][0] ), .C(
        \ImageBuffer[38][0] ), .D(\ImageBuffer[39][0] ), .S0(n4114), .S1(n4131), .Y(n3956) );
  MX4X1 U6406 ( .A(\ImageBuffer[36][2] ), .B(\ImageBuffer[37][2] ), .C(
        \ImageBuffer[38][2] ), .D(\ImageBuffer[39][2] ), .S0(n3939), .S1(n3930), .Y(n3807) );
  MX4X1 U6407 ( .A(\ImageBuffer[4][2] ), .B(\ImageBuffer[5][2] ), .C(
        \ImageBuffer[6][2] ), .D(\ImageBuffer[7][2] ), .S0(n3939), .S1(n3926), 
        .Y(n3817) );
  MX4X1 U6408 ( .A(\ImageBuffer[52][0] ), .B(\ImageBuffer[53][0] ), .C(
        \ImageBuffer[54][0] ), .D(\ImageBuffer[55][0] ), .S0(n4117), .S1(n3749), .Y(n3575) );
  MX4X1 U6409 ( .A(\ImageBuffer[36][0] ), .B(\ImageBuffer[37][0] ), .C(
        \ImageBuffer[38][0] ), .D(\ImageBuffer[39][0] ), .S0(n4117), .S1(n3750), .Y(n3580) );
  MX4X1 U6410 ( .A(\ImageBuffer[20][0] ), .B(\ImageBuffer[21][0] ), .C(
        \ImageBuffer[22][0] ), .D(\ImageBuffer[23][0] ), .S0(n3512), .S1(n3473), .Y(n4331) );
  MX4X1 U6411 ( .A(\ImageBuffer[52][0] ), .B(\ImageBuffer[53][0] ), .C(
        \ImageBuffer[54][0] ), .D(\ImageBuffer[55][0] ), .S0(n3938), .S1(n3923), .Y(n3762) );
  MX4X1 U6412 ( .A(\ImageBuffer[36][0] ), .B(\ImageBuffer[37][0] ), .C(
        \ImageBuffer[38][0] ), .D(\ImageBuffer[39][0] ), .S0(n3938), .S1(n3920), .Y(n3767) );
  MX4X1 U6413 ( .A(\ImageBuffer[20][2] ), .B(\ImageBuffer[21][2] ), .C(
        \ImageBuffer[22][2] ), .D(\ImageBuffer[23][2] ), .S0(n3740), .S1(n4132), .Y(n4000) );
  MX4X1 U6414 ( .A(\ImageBuffer[52][2] ), .B(\ImageBuffer[53][2] ), .C(
        \ImageBuffer[54][2] ), .D(\ImageBuffer[55][2] ), .S0(n4115), .S1(n3749), .Y(n3990) );
  MX4X1 U6415 ( .A(\ImageBuffer[4][0] ), .B(\ImageBuffer[5][0] ), .C(
        \ImageBuffer[6][0] ), .D(\ImageBuffer[7][0] ), .S0(n3740), .S1(n4128), 
        .Y(n3590) );
  MX4X1 U6416 ( .A(\ImageBuffer[20][2] ), .B(\ImageBuffer[21][2] ), .C(
        \ImageBuffer[22][2] ), .D(\ImageBuffer[23][2] ), .S0(n3939), .S1(n5123), .Y(n3812) );
  MX4X1 U6417 ( .A(\ImageBuffer[52][2] ), .B(\ImageBuffer[53][2] ), .C(
        \ImageBuffer[54][2] ), .D(\ImageBuffer[55][2] ), .S0(n5120), .S1(n3927), .Y(n3802) );
  MX4X1 U6418 ( .A(\ImageBuffer[4][0] ), .B(\ImageBuffer[5][0] ), .C(
        \ImageBuffer[6][0] ), .D(\ImageBuffer[7][0] ), .S0(n3939), .S1(n3922), 
        .Y(n3777) );
  MX4X1 U6419 ( .A(\ImageBuffer[52][0] ), .B(\ImageBuffer[53][0] ), .C(
        \ImageBuffer[54][0] ), .D(\ImageBuffer[55][0] ), .S0(n3519), .S1(n3472), .Y(n4321) );
  MX4X1 U6420 ( .A(\ImageBuffer[52][2] ), .B(\ImageBuffer[53][2] ), .C(
        \ImageBuffer[54][2] ), .D(\ImageBuffer[55][2] ), .S0(n3347), .S1(n3482), .Y(n4521) );
  MX4X1 U6421 ( .A(\ImageBuffer[4][2] ), .B(\ImageBuffer[5][2] ), .C(
        \ImageBuffer[6][2] ), .D(\ImageBuffer[7][2] ), .S0(n3506), .S1(n3483), 
        .Y(n4536) );
  MX4X1 U6422 ( .A(\ImageBuffer[20][2] ), .B(\ImageBuffer[21][2] ), .C(
        \ImageBuffer[22][2] ), .D(\ImageBuffer[23][2] ), .S0(n3741), .S1(n3752), .Y(n3625) );
  MX4X1 U6423 ( .A(\ImageBuffer[52][2] ), .B(\ImageBuffer[53][2] ), .C(
        \ImageBuffer[54][2] ), .D(\ImageBuffer[55][2] ), .S0(n4119), .S1(n4124), .Y(n3615) );
  MX4X1 U6424 ( .A(\ImageBuffer[36][2] ), .B(\ImageBuffer[37][2] ), .C(
        \ImageBuffer[38][2] ), .D(\ImageBuffer[39][2] ), .S0(n3741), .S1(n3751), .Y(n3620) );
  MX4X1 U6425 ( .A(\ImageBuffer[4][2] ), .B(\ImageBuffer[5][2] ), .C(
        \ImageBuffer[6][2] ), .D(\ImageBuffer[7][2] ), .S0(n3741), .S1(N2494), 
        .Y(n3630) );
  MX4X1 U6426 ( .A(\ImageBuffer[20][3] ), .B(\ImageBuffer[21][3] ), .C(
        \ImageBuffer[22][3] ), .D(\ImageBuffer[23][3] ), .S0(n3498), .S1(n4122), .Y(n3645) );
  MX4X1 U6427 ( .A(\ImageBuffer[52][3] ), .B(\ImageBuffer[53][3] ), .C(
        \ImageBuffer[54][3] ), .D(\ImageBuffer[55][3] ), .S0(n3498), .S1(n4128), .Y(n3635) );
  MX4X1 U6428 ( .A(\ImageBuffer[36][3] ), .B(\ImageBuffer[37][3] ), .C(
        \ImageBuffer[38][3] ), .D(\ImageBuffer[39][3] ), .S0(n3498), .S1(n3756), .Y(n3640) );
  MX4X1 U6429 ( .A(\ImageBuffer[4][3] ), .B(\ImageBuffer[5][3] ), .C(
        \ImageBuffer[6][3] ), .D(\ImageBuffer[7][3] ), .S0(n3498), .S1(n4129), 
        .Y(n3650) );
  MX4X1 U6430 ( .A(\ImageBuffer[20][6] ), .B(\ImageBuffer[21][6] ), .C(
        \ImageBuffer[22][6] ), .D(\ImageBuffer[23][6] ), .S0(n3488), .S1(n3756), .Y(n3705) );
  MX4X1 U6431 ( .A(\ImageBuffer[52][6] ), .B(\ImageBuffer[53][6] ), .C(
        \ImageBuffer[54][6] ), .D(\ImageBuffer[55][6] ), .S0(n3743), .S1(n4128), .Y(n3695) );
  MX4X1 U6432 ( .A(\ImageBuffer[20][5] ), .B(\ImageBuffer[21][5] ), .C(
        \ImageBuffer[22][5] ), .D(\ImageBuffer[23][5] ), .S0(n4117), .S1(n4131), .Y(n4060) );
  MX4X1 U6433 ( .A(\ImageBuffer[4][5] ), .B(\ImageBuffer[5][5] ), .C(
        \ImageBuffer[6][5] ), .D(\ImageBuffer[7][5] ), .S0(n4117), .S1(n4125), 
        .Y(n4065) );
  MX4X1 U6434 ( .A(\ImageBuffer[52][6] ), .B(\ImageBuffer[53][6] ), .C(
        \ImageBuffer[54][6] ), .D(\ImageBuffer[55][6] ), .S0(n4117), .S1(n4131), .Y(n4070) );
  MX4X1 U6435 ( .A(\ImageBuffer[52][3] ), .B(\ImageBuffer[53][3] ), .C(
        \ImageBuffer[54][3] ), .D(\ImageBuffer[55][3] ), .S0(n4116), .S1(n4125), .Y(n4010) );
  MX4X1 U6436 ( .A(\ImageBuffer[4][3] ), .B(\ImageBuffer[5][3] ), .C(
        \ImageBuffer[6][3] ), .D(\ImageBuffer[7][3] ), .S0(n4116), .S1(n4130), 
        .Y(n4025) );
  MX4X1 U6437 ( .A(\ImageBuffer[52][3] ), .B(\ImageBuffer[53][3] ), .C(
        \ImageBuffer[54][3] ), .D(\ImageBuffer[55][3] ), .S0(n3489), .S1(n3927), .Y(n3822) );
  MX4X1 U6438 ( .A(\ImageBuffer[36][3] ), .B(\ImageBuffer[37][3] ), .C(
        \ImageBuffer[38][3] ), .D(\ImageBuffer[39][3] ), .S0(n3489), .S1(n3920), .Y(n3827) );
  MX4X1 U6439 ( .A(\ImageBuffer[52][4] ), .B(\ImageBuffer[53][4] ), .C(
        \ImageBuffer[54][4] ), .D(\ImageBuffer[55][4] ), .S0(n3742), .S1(n4127), .Y(n3655) );
  MX4X1 U6440 ( .A(\ImageBuffer[4][4] ), .B(\ImageBuffer[5][4] ), .C(
        \ImageBuffer[6][4] ), .D(\ImageBuffer[7][4] ), .S0(n3498), .S1(n4128), 
        .Y(n3670) );
  MX4X1 U6441 ( .A(\ImageBuffer[36][4] ), .B(\ImageBuffer[37][4] ), .C(
        \ImageBuffer[38][4] ), .D(\ImageBuffer[39][4] ), .S0(n3486), .S1(n3927), .Y(n3847) );
  MX4X1 U6442 ( .A(\ImageBuffer[4][4] ), .B(\ImageBuffer[5][4] ), .C(
        \ImageBuffer[6][4] ), .D(\ImageBuffer[7][4] ), .S0(n3941), .S1(n3920), 
        .Y(n3857) );
  MX4X1 U6443 ( .A(\ImageBuffer[20][1] ), .B(\ImageBuffer[21][1] ), .C(
        \ImageBuffer[22][1] ), .D(\ImageBuffer[23][1] ), .S0(n3736), .S1(n4134), .Y(n3605) );
  MX4X1 U6444 ( .A(\ImageBuffer[20][2] ), .B(\ImageBuffer[21][2] ), .C(
        \ImageBuffer[22][2] ), .D(\ImageBuffer[23][2] ), .S0(n3938), .S1(n4311), .Y(n4189) );
  MX4X1 U6445 ( .A(\ImageBuffer[52][2] ), .B(\ImageBuffer[53][2] ), .C(
        \ImageBuffer[54][2] ), .D(\ImageBuffer[55][2] ), .S0(n4300), .S1(n4311), .Y(n4179) );
  MX4X1 U6446 ( .A(\ImageBuffer[4][2] ), .B(\ImageBuffer[5][2] ), .C(
        \ImageBuffer[6][2] ), .D(\ImageBuffer[7][2] ), .S0(n3938), .S1(n4312), 
        .Y(n4194) );
  MX4X1 U6447 ( .A(\ImageBuffer[36][2] ), .B(\ImageBuffer[37][2] ), .C(
        \ImageBuffer[38][2] ), .D(\ImageBuffer[39][2] ), .S0(n3938), .S1(n4306), .Y(n4184) );
  MX4X1 U6448 ( .A(\ImageBuffer[20][6] ), .B(\ImageBuffer[21][6] ), .C(
        \ImageBuffer[22][6] ), .D(\ImageBuffer[23][6] ), .S0(n3939), .S1(n3925), .Y(n3892) );
  MX4X1 U6449 ( .A(\ImageBuffer[36][6] ), .B(\ImageBuffer[37][6] ), .C(
        \ImageBuffer[38][6] ), .D(\ImageBuffer[39][6] ), .S0(n3939), .S1(n3920), .Y(n3887) );
  MX4X1 U6450 ( .A(\ImageBuffer[4][6] ), .B(\ImageBuffer[5][6] ), .C(
        \ImageBuffer[6][6] ), .D(\ImageBuffer[7][6] ), .S0(n3939), .S1(n3931), 
        .Y(n3897) );
  MX4X1 U6451 ( .A(\ImageBuffer[36][4] ), .B(\ImageBuffer[37][4] ), .C(
        \ImageBuffer[38][4] ), .D(\ImageBuffer[39][4] ), .S0(n4300), .S1(n4312), .Y(n4224) );
  MX4X1 U6452 ( .A(\ImageBuffer[20][4] ), .B(\ImageBuffer[21][4] ), .C(
        \ImageBuffer[22][4] ), .D(\ImageBuffer[23][4] ), .S0(n3486), .S1(n4310), .Y(n4229) );
  MX4X1 U6453 ( .A(\ImageBuffer[52][4] ), .B(\ImageBuffer[53][4] ), .C(
        \ImageBuffer[54][4] ), .D(\ImageBuffer[55][4] ), .S0(n3941), .S1(n4308), .Y(n4219) );
  MX4X1 U6454 ( .A(\ImageBuffer[20][6] ), .B(\ImageBuffer[21][6] ), .C(
        \ImageBuffer[22][6] ), .D(\ImageBuffer[23][6] ), .S0(n4297), .S1(n4311), .Y(n4269) );
  MX4X1 U6455 ( .A(\ImageBuffer[4][6] ), .B(\ImageBuffer[5][6] ), .C(
        \ImageBuffer[6][6] ), .D(\ImageBuffer[7][6] ), .S0(n4300), .S1(n4313), 
        .Y(n4274) );
  MX4X1 U6456 ( .A(\ImageBuffer[36][6] ), .B(\ImageBuffer[37][6] ), .C(
        \ImageBuffer[38][6] ), .D(\ImageBuffer[39][6] ), .S0(n4300), .S1(n4314), .Y(n4264) );
  MX4X1 U6457 ( .A(\ImageBuffer[52][0] ), .B(\ImageBuffer[53][0] ), .C(
        \ImageBuffer[54][0] ), .D(\ImageBuffer[55][0] ), .S0(n3938), .S1(n4310), .Y(n4139) );
  MX4X1 U6458 ( .A(\ImageBuffer[4][0] ), .B(\ImageBuffer[5][0] ), .C(
        \ImageBuffer[6][0] ), .D(\ImageBuffer[7][0] ), .S0(n3939), .S1(n4316), 
        .Y(n4154) );
  MX4X1 U6459 ( .A(\ImageBuffer[36][0] ), .B(\ImageBuffer[37][0] ), .C(
        \ImageBuffer[38][0] ), .D(\ImageBuffer[39][0] ), .S0(n3938), .S1(n4308), .Y(n4144) );
  MX4X1 U6460 ( .A(\ImageBuffer[4][0] ), .B(\ImageBuffer[5][0] ), .C(
        \ImageBuffer[6][0] ), .D(\ImageBuffer[7][0] ), .S0(n3521), .S1(n3474), 
        .Y(n4336) );
  MX4X1 U6461 ( .A(\ImageBuffer[36][0] ), .B(\ImageBuffer[37][0] ), .C(
        \ImageBuffer[38][0] ), .D(\ImageBuffer[39][0] ), .S0(n3519), .S1(n3473), .Y(n4326) );
  MX4X1 U6462 ( .A(\ImageBuffer[4][0] ), .B(\ImageBuffer[5][0] ), .C(
        \ImageBuffer[6][0] ), .D(\ImageBuffer[7][0] ), .S0(n3343), .S1(n3483), 
        .Y(n4496) );
  MX4X1 U6463 ( .A(\ImageBuffer[52][0] ), .B(\ImageBuffer[53][0] ), .C(
        \ImageBuffer[54][0] ), .D(\ImageBuffer[55][0] ), .S0(n3347), .S1(n3483), .Y(n4481) );
  MX4X1 U6464 ( .A(\ImageBuffer[36][0] ), .B(\ImageBuffer[37][0] ), .C(
        \ImageBuffer[38][0] ), .D(\ImageBuffer[39][0] ), .S0(n3343), .S1(n3482), .Y(n4486) );
  MX4X1 U6465 ( .A(\ImageBuffer[52][1] ), .B(\ImageBuffer[53][1] ), .C(
        \ImageBuffer[54][1] ), .D(\ImageBuffer[55][1] ), .S0(n3506), .S1(n3484), .Y(n4501) );
  MX4X1 U6466 ( .A(\ImageBuffer[20][1] ), .B(\ImageBuffer[21][1] ), .C(
        \ImageBuffer[22][1] ), .D(\ImageBuffer[23][1] ), .S0(n3343), .S1(n3482), .Y(n4511) );
  MX4X1 U6467 ( .A(\ImageBuffer[36][1] ), .B(\ImageBuffer[37][1] ), .C(
        \ImageBuffer[38][1] ), .D(\ImageBuffer[39][1] ), .S0(n3343), .S1(n3482), .Y(n4506) );
  MX4X1 U6468 ( .A(\ImageBuffer[4][1] ), .B(\ImageBuffer[5][1] ), .C(
        \ImageBuffer[6][1] ), .D(\ImageBuffer[7][1] ), .S0(n3347), .S1(n3482), 
        .Y(n4516) );
  MX4X1 U6469 ( .A(\ImageBuffer[36][1] ), .B(\ImageBuffer[37][1] ), .C(
        \ImageBuffer[38][1] ), .D(\ImageBuffer[39][1] ), .S0(n3513), .S1(n3473), .Y(n4346) );
  MX4X1 U6470 ( .A(\ImageBuffer[4][1] ), .B(\ImageBuffer[5][1] ), .C(
        \ImageBuffer[6][1] ), .D(\ImageBuffer[7][1] ), .S0(n3515), .S1(n3472), 
        .Y(n4356) );
  MX4X1 U6471 ( .A(\ImageBuffer[36][3] ), .B(\ImageBuffer[37][3] ), .C(
        \ImageBuffer[38][3] ), .D(\ImageBuffer[39][3] ), .S0(n3522), .S1(n3472), .Y(n4386) );
  MX4X1 U6472 ( .A(\ImageBuffer[4][3] ), .B(\ImageBuffer[5][3] ), .C(
        \ImageBuffer[6][3] ), .D(\ImageBuffer[7][3] ), .S0(n3511), .S1(n3471), 
        .Y(n4396) );
  MX4X1 U6473 ( .A(\ImageBuffer[20][3] ), .B(\ImageBuffer[21][3] ), .C(
        \ImageBuffer[22][3] ), .D(\ImageBuffer[23][3] ), .S0(n3506), .S1(n3484), .Y(n4551) );
  MX4X1 U6474 ( .A(\ImageBuffer[36][3] ), .B(\ImageBuffer[37][3] ), .C(
        \ImageBuffer[38][3] ), .D(\ImageBuffer[39][3] ), .S0(n3343), .S1(n3485), .Y(n4546) );
  MX4X1 U6475 ( .A(\ImageBuffer[4][3] ), .B(\ImageBuffer[5][3] ), .C(
        \ImageBuffer[6][3] ), .D(\ImageBuffer[7][3] ), .S0(n3347), .S1(n3482), 
        .Y(n4556) );
  MX4X1 U6476 ( .A(\ImageBuffer[20][4] ), .B(\ImageBuffer[21][4] ), .C(
        \ImageBuffer[22][4] ), .D(\ImageBuffer[23][4] ), .S0(n3514), .S1(n3473), .Y(n4411) );
  MX4X1 U6477 ( .A(\ImageBuffer[52][4] ), .B(\ImageBuffer[53][4] ), .C(
        \ImageBuffer[54][4] ), .D(\ImageBuffer[55][4] ), .S0(n3511), .S1(n3471), .Y(n4401) );
  MX4X1 U6478 ( .A(\ImageBuffer[36][4] ), .B(\ImageBuffer[37][4] ), .C(
        \ImageBuffer[38][4] ), .D(\ImageBuffer[39][4] ), .S0(n3517), .S1(n3473), .Y(n4406) );
  MX4X1 U6479 ( .A(\ImageBuffer[4][4] ), .B(\ImageBuffer[5][4] ), .C(
        \ImageBuffer[6][4] ), .D(\ImageBuffer[7][4] ), .S0(n3513), .S1(n3471), 
        .Y(n4416) );
  MX4X1 U6480 ( .A(\ImageBuffer[20][4] ), .B(\ImageBuffer[21][4] ), .C(
        \ImageBuffer[22][4] ), .D(\ImageBuffer[23][4] ), .S0(n3506), .S1(n3484), .Y(n4571) );
  MX4X1 U6481 ( .A(\ImageBuffer[52][4] ), .B(\ImageBuffer[53][4] ), .C(
        \ImageBuffer[54][4] ), .D(\ImageBuffer[55][4] ), .S0(n3347), .S1(n3485), .Y(n4561) );
  MX4X1 U6482 ( .A(\ImageBuffer[36][4] ), .B(\ImageBuffer[37][4] ), .C(
        \ImageBuffer[38][4] ), .D(\ImageBuffer[39][4] ), .S0(n3343), .S1(n3485), .Y(n4566) );
  MX4X1 U6483 ( .A(\ImageBuffer[4][4] ), .B(\ImageBuffer[5][4] ), .C(
        \ImageBuffer[6][4] ), .D(\ImageBuffer[7][4] ), .S0(n3347), .S1(n3482), 
        .Y(n4576) );
  MX4X1 U6484 ( .A(\ImageBuffer[20][5] ), .B(\ImageBuffer[21][5] ), .C(
        \ImageBuffer[22][5] ), .D(\ImageBuffer[23][5] ), .S0(n3515), .S1(n3473), .Y(n4431) );
  MX4X1 U6485 ( .A(\ImageBuffer[52][5] ), .B(\ImageBuffer[53][5] ), .C(
        \ImageBuffer[54][5] ), .D(\ImageBuffer[55][5] ), .S0(n3522), .S1(n3471), .Y(n4421) );
  MX4X1 U6486 ( .A(\ImageBuffer[36][5] ), .B(\ImageBuffer[37][5] ), .C(
        \ImageBuffer[38][5] ), .D(\ImageBuffer[39][5] ), .S0(n3511), .S1(n3472), .Y(n4426) );
  MX4X1 U6487 ( .A(\ImageBuffer[4][5] ), .B(\ImageBuffer[5][5] ), .C(
        \ImageBuffer[6][5] ), .D(\ImageBuffer[7][5] ), .S0(n3516), .S1(n3471), 
        .Y(n4436) );
  MX4X1 U6488 ( .A(\ImageBuffer[20][5] ), .B(\ImageBuffer[21][5] ), .C(
        \ImageBuffer[22][5] ), .D(\ImageBuffer[23][5] ), .S0(n3343), .S1(n3484), .Y(n4591) );
  MX4X1 U6489 ( .A(\ImageBuffer[52][5] ), .B(\ImageBuffer[53][5] ), .C(
        \ImageBuffer[54][5] ), .D(\ImageBuffer[55][5] ), .S0(n3343), .S1(n3483), .Y(n4581) );
  MX4X1 U6490 ( .A(\ImageBuffer[36][5] ), .B(\ImageBuffer[37][5] ), .C(
        \ImageBuffer[38][5] ), .D(\ImageBuffer[39][5] ), .S0(n3347), .S1(n3484), .Y(n4586) );
  MX4X1 U6491 ( .A(\ImageBuffer[4][5] ), .B(\ImageBuffer[5][5] ), .C(
        \ImageBuffer[6][5] ), .D(\ImageBuffer[7][5] ), .S0(n3506), .S1(n3485), 
        .Y(n4596) );
  MX4X1 U6492 ( .A(\ImageBuffer[20][6] ), .B(\ImageBuffer[21][6] ), .C(
        \ImageBuffer[22][6] ), .D(\ImageBuffer[23][6] ), .S0(n3521), .S1(n3473), .Y(n4451) );
  MX4X1 U6493 ( .A(\ImageBuffer[52][6] ), .B(\ImageBuffer[53][6] ), .C(
        \ImageBuffer[54][6] ), .D(\ImageBuffer[55][6] ), .S0(n3512), .S1(n3472), .Y(n4441) );
  MX4X1 U6494 ( .A(\ImageBuffer[36][6] ), .B(\ImageBuffer[37][6] ), .C(
        \ImageBuffer[38][6] ), .D(\ImageBuffer[39][6] ), .S0(n3511), .S1(n3474), .Y(n4446) );
  MX4X1 U6495 ( .A(\ImageBuffer[4][6] ), .B(\ImageBuffer[5][6] ), .C(
        \ImageBuffer[6][6] ), .D(\ImageBuffer[7][6] ), .S0(n3514), .S1(n3473), 
        .Y(n4456) );
  MX4X1 U6496 ( .A(\ImageBuffer[20][6] ), .B(\ImageBuffer[21][6] ), .C(
        \ImageBuffer[22][6] ), .D(\ImageBuffer[23][6] ), .S0(n3347), .S1(n3485), .Y(n4611) );
  MX4X1 U6497 ( .A(\ImageBuffer[52][6] ), .B(\ImageBuffer[53][6] ), .C(
        \ImageBuffer[54][6] ), .D(\ImageBuffer[55][6] ), .S0(n3343), .S1(n3484), .Y(n4601) );
  MX4X1 U6498 ( .A(\ImageBuffer[36][6] ), .B(\ImageBuffer[37][6] ), .C(
        \ImageBuffer[38][6] ), .D(\ImageBuffer[39][6] ), .S0(n3347), .S1(n3482), .Y(n4606) );
  MX4X1 U6499 ( .A(\ImageBuffer[4][6] ), .B(\ImageBuffer[5][6] ), .C(
        \ImageBuffer[6][6] ), .D(\ImageBuffer[7][6] ), .S0(n3347), .S1(n3484), 
        .Y(n4616) );
  MX4X1 U6500 ( .A(\ImageBuffer[20][7] ), .B(\ImageBuffer[21][7] ), .C(
        \ImageBuffer[22][7] ), .D(\ImageBuffer[23][7] ), .S0(n3513), .S1(n3473), .Y(n4471) );
  MX4X1 U6501 ( .A(\ImageBuffer[52][7] ), .B(\ImageBuffer[53][7] ), .C(
        \ImageBuffer[54][7] ), .D(\ImageBuffer[55][7] ), .S0(n3516), .S1(n3473), .Y(n4461) );
  MX4X1 U6502 ( .A(\ImageBuffer[36][7] ), .B(\ImageBuffer[37][7] ), .C(
        \ImageBuffer[38][7] ), .D(\ImageBuffer[39][7] ), .S0(n3522), .S1(n3474), .Y(n4466) );
  MX4X1 U6503 ( .A(\ImageBuffer[4][7] ), .B(\ImageBuffer[5][7] ), .C(
        \ImageBuffer[6][7] ), .D(\ImageBuffer[7][7] ), .S0(n3513), .S1(n3471), 
        .Y(n4476) );
  MX4X1 U6504 ( .A(\ImageBuffer[20][7] ), .B(\ImageBuffer[21][7] ), .C(
        \ImageBuffer[22][7] ), .D(\ImageBuffer[23][7] ), .S0(n3506), .S1(n3484), .Y(n4631) );
  MX4X1 U6505 ( .A(\ImageBuffer[52][7] ), .B(\ImageBuffer[53][7] ), .C(
        \ImageBuffer[54][7] ), .D(\ImageBuffer[55][7] ), .S0(n3346), .S1(n3483), .Y(n4621) );
  MX4X1 U6506 ( .A(\ImageBuffer[36][7] ), .B(\ImageBuffer[37][7] ), .C(
        \ImageBuffer[38][7] ), .D(\ImageBuffer[39][7] ), .S0(n3342), .S1(n3485), .Y(n4626) );
  MX4X1 U6507 ( .A(\ImageBuffer[4][7] ), .B(\ImageBuffer[5][7] ), .C(
        \ImageBuffer[6][7] ), .D(\ImageBuffer[7][7] ), .S0(n3346), .S1(n3483), 
        .Y(n4636) );
  MX4X1 U6508 ( .A(\ImageBuffer[20][4] ), .B(\ImageBuffer[21][4] ), .C(
        \ImageBuffer[22][4] ), .D(\ImageBuffer[23][4] ), .S0(n4119), .S1(n4125), .Y(n4040) );
  MX4X1 U6509 ( .A(\ImageBuffer[52][4] ), .B(\ImageBuffer[53][4] ), .C(
        \ImageBuffer[54][4] ), .D(\ImageBuffer[55][4] ), .S0(n4119), .S1(n4127), .Y(n4030) );
  MX4X1 U6510 ( .A(\ImageBuffer[36][4] ), .B(\ImageBuffer[37][4] ), .C(
        \ImageBuffer[38][4] ), .D(\ImageBuffer[39][4] ), .S0(n4119), .S1(n3750), .Y(n4035) );
  MX4X1 U6511 ( .A(\ImageBuffer[4][4] ), .B(\ImageBuffer[5][4] ), .C(
        \ImageBuffer[6][4] ), .D(\ImageBuffer[7][4] ), .S0(n3737), .S1(n4134), 
        .Y(n4045) );
  MX4X1 U6512 ( .A(\ImageBuffer[24][0] ), .B(\ImageBuffer[25][0] ), .C(
        \ImageBuffer[26][0] ), .D(\ImageBuffer[27][0] ), .S0(n3939), .S1(n4311), .Y(n4148) );
  MX4X1 U6513 ( .A(\ImageBuffer[28][0] ), .B(\ImageBuffer[29][0] ), .C(
        \ImageBuffer[30][0] ), .D(\ImageBuffer[31][0] ), .S0(n3938), .S1(n4315), .Y(n4147) );
  MX4X1 U6514 ( .A(\ImageBuffer[20][0] ), .B(\ImageBuffer[21][0] ), .C(
        \ImageBuffer[22][0] ), .D(\ImageBuffer[23][0] ), .S0(n3939), .S1(n4316), .Y(n4149) );
  MX4X1 U6515 ( .A(\ImageBuffer[16][2] ), .B(\ImageBuffer[17][2] ), .C(
        \ImageBuffer[18][2] ), .D(\ImageBuffer[19][2] ), .S0(n3740), .S1(n4126), .Y(n4001) );
  MX4X1 U6516 ( .A(\ImageBuffer[24][2] ), .B(\ImageBuffer[25][2] ), .C(
        \ImageBuffer[26][2] ), .D(\ImageBuffer[27][2] ), .S0(n3740), .S1(n4129), .Y(n3999) );
  MX4X1 U6517 ( .A(\ImageBuffer[28][2] ), .B(\ImageBuffer[29][2] ), .C(
        \ImageBuffer[30][2] ), .D(\ImageBuffer[31][2] ), .S0(n3735), .S1(n4124), .Y(n3998) );
  MX4X1 U6518 ( .A(\ImageBuffer[16][6] ), .B(\ImageBuffer[17][6] ), .C(
        \ImageBuffer[18][6] ), .D(\ImageBuffer[19][6] ), .S0(n3939), .S1(n3499), .Y(n3893) );
  MX4X1 U6519 ( .A(\ImageBuffer[24][6] ), .B(\ImageBuffer[25][6] ), .C(
        \ImageBuffer[26][6] ), .D(\ImageBuffer[27][6] ), .S0(n4297), .S1(n3925), .Y(n3891) );
  MX4X1 U6520 ( .A(\ImageBuffer[28][6] ), .B(\ImageBuffer[29][6] ), .C(
        \ImageBuffer[30][6] ), .D(\ImageBuffer[31][6] ), .S0(n4297), .S1(n3923), .Y(n3890) );
  MX4X1 U6521 ( .A(\ImageBuffer[16][4] ), .B(\ImageBuffer[17][4] ), .C(
        \ImageBuffer[18][4] ), .D(\ImageBuffer[19][4] ), .S0(n3506), .S1(n3484), .Y(n4572) );
  MX4X1 U6522 ( .A(\ImageBuffer[24][4] ), .B(\ImageBuffer[25][4] ), .C(
        \ImageBuffer[26][4] ), .D(\ImageBuffer[27][4] ), .S0(n3506), .S1(n3484), .Y(n4570) );
  MX4X1 U6523 ( .A(\ImageBuffer[28][4] ), .B(\ImageBuffer[29][4] ), .C(
        \ImageBuffer[30][4] ), .D(\ImageBuffer[31][4] ), .S0(n3343), .S1(n3482), .Y(n4569) );
  MX4X1 U6524 ( .A(n4592), .B(n4590), .C(n4591), .D(n4589), .S0(n3496), .S1(
        n4640), .Y(n4593) );
  MX4X1 U6525 ( .A(\ImageBuffer[16][5] ), .B(\ImageBuffer[17][5] ), .C(
        \ImageBuffer[18][5] ), .D(\ImageBuffer[19][5] ), .S0(n3506), .S1(n3483), .Y(n4592) );
  MX4X1 U6526 ( .A(\ImageBuffer[24][5] ), .B(\ImageBuffer[25][5] ), .C(
        \ImageBuffer[26][5] ), .D(\ImageBuffer[27][5] ), .S0(n3343), .S1(n3483), .Y(n4590) );
  MX4X1 U6527 ( .A(\ImageBuffer[28][5] ), .B(\ImageBuffer[29][5] ), .C(
        \ImageBuffer[30][5] ), .D(\ImageBuffer[31][5] ), .S0(n3506), .S1(n3482), .Y(n4589) );
  MX4X1 U6528 ( .A(n4452), .B(n4450), .C(n4451), .D(n4449), .S0(n3503), .S1(
        n3495), .Y(n4453) );
  MX4X1 U6529 ( .A(\ImageBuffer[16][6] ), .B(\ImageBuffer[17][6] ), .C(
        \ImageBuffer[18][6] ), .D(\ImageBuffer[19][6] ), .S0(n3513), .S1(n3473), .Y(n4452) );
  MX4X1 U6530 ( .A(\ImageBuffer[24][6] ), .B(\ImageBuffer[25][6] ), .C(
        \ImageBuffer[26][6] ), .D(\ImageBuffer[27][6] ), .S0(n3522), .S1(n3471), .Y(n4450) );
  MX4X1 U6531 ( .A(\ImageBuffer[28][6] ), .B(\ImageBuffer[29][6] ), .C(
        \ImageBuffer[30][6] ), .D(\ImageBuffer[31][6] ), .S0(n3519), .S1(n3471), .Y(n4449) );
  MX4X1 U6532 ( .A(\ImageBuffer[16][2] ), .B(\ImageBuffer[17][2] ), .C(
        \ImageBuffer[18][2] ), .D(\ImageBuffer[19][2] ), .S0(n3938), .S1(n4303), .Y(n4190) );
  MX4X1 U6533 ( .A(\ImageBuffer[24][2] ), .B(\ImageBuffer[25][2] ), .C(
        \ImageBuffer[26][2] ), .D(\ImageBuffer[27][2] ), .S0(n3938), .S1(n4312), .Y(n4188) );
  MX4X1 U6534 ( .A(\ImageBuffer[28][2] ), .B(\ImageBuffer[29][2] ), .C(
        \ImageBuffer[30][2] ), .D(\ImageBuffer[31][2] ), .S0(n3938), .S1(n4307), .Y(n4187) );
  MX4X1 U6535 ( .A(\ImageBuffer[32][2] ), .B(\ImageBuffer[33][2] ), .C(
        \ImageBuffer[34][2] ), .D(\ImageBuffer[35][2] ), .S0(n3740), .S1(n3755), .Y(n3996) );
  MX4X1 U6536 ( .A(\ImageBuffer[0][2] ), .B(\ImageBuffer[1][2] ), .C(
        \ImageBuffer[2][2] ), .D(\ImageBuffer[3][2] ), .S0(n3740), .S1(n3749), 
        .Y(n4006) );
  MX4X1 U6537 ( .A(\ImageBuffer[48][0] ), .B(\ImageBuffer[49][0] ), .C(
        \ImageBuffer[50][0] ), .D(\ImageBuffer[51][0] ), .S0(n4114), .S1(n4131), .Y(n3953) );
  MX4X1 U6538 ( .A(\ImageBuffer[32][2] ), .B(\ImageBuffer[33][2] ), .C(
        \ImageBuffer[34][2] ), .D(\ImageBuffer[35][2] ), .S0(n3939), .S1(n3931), .Y(n3808) );
  MX4X1 U6539 ( .A(\ImageBuffer[0][2] ), .B(\ImageBuffer[1][2] ), .C(
        \ImageBuffer[2][2] ), .D(\ImageBuffer[3][2] ), .S0(n3939), .S1(n3341), 
        .Y(n3818) );
  MX4X1 U6540 ( .A(\ImageBuffer[48][0] ), .B(\ImageBuffer[49][0] ), .C(
        \ImageBuffer[50][0] ), .D(\ImageBuffer[51][0] ), .S0(n4117), .S1(n3756), .Y(n3576) );
  MX4X1 U6541 ( .A(\ImageBuffer[32][0] ), .B(\ImageBuffer[33][0] ), .C(
        \ImageBuffer[34][0] ), .D(\ImageBuffer[35][0] ), .S0(n4119), .S1(n3748), .Y(n3581) );
  MX4X1 U6542 ( .A(\ImageBuffer[16][0] ), .B(\ImageBuffer[17][0] ), .C(
        \ImageBuffer[18][0] ), .D(\ImageBuffer[19][0] ), .S0(n3519), .S1(n3472), .Y(n4332) );
  MX4X1 U6543 ( .A(\ImageBuffer[48][0] ), .B(\ImageBuffer[49][0] ), .C(
        \ImageBuffer[50][0] ), .D(\ImageBuffer[51][0] ), .S0(n3938), .S1(n3920), .Y(n3763) );
  MX4X1 U6544 ( .A(\ImageBuffer[32][0] ), .B(\ImageBuffer[33][0] ), .C(
        \ImageBuffer[34][0] ), .D(\ImageBuffer[35][0] ), .S0(n3938), .S1(n3923), .Y(n3768) );
  MX4X1 U6545 ( .A(\ImageBuffer[16][0] ), .B(\ImageBuffer[17][0] ), .C(
        \ImageBuffer[18][0] ), .D(\ImageBuffer[19][0] ), .S0(n3939), .S1(n3480), .Y(n3773) );
  MX4X1 U6546 ( .A(\ImageBuffer[48][2] ), .B(\ImageBuffer[49][2] ), .C(
        \ImageBuffer[50][2] ), .D(\ImageBuffer[51][2] ), .S0(n3343), .S1(n3484), .Y(n4522) );
  MX4X1 U6547 ( .A(\ImageBuffer[0][2] ), .B(\ImageBuffer[1][2] ), .C(
        \ImageBuffer[2][2] ), .D(\ImageBuffer[3][2] ), .S0(n3347), .S1(n3484), 
        .Y(n4537) );
  MX4X1 U6548 ( .A(\ImageBuffer[32][2] ), .B(\ImageBuffer[33][2] ), .C(
        \ImageBuffer[34][2] ), .D(\ImageBuffer[35][2] ), .S0(n3741), .S1(n4129), .Y(n3621) );
  MX4X1 U6549 ( .A(\ImageBuffer[0][2] ), .B(\ImageBuffer[1][2] ), .C(
        \ImageBuffer[2][2] ), .D(\ImageBuffer[3][2] ), .S0(n3741), .S1(n3753), 
        .Y(n3631) );
  MX4X1 U6550 ( .A(\ImageBuffer[32][3] ), .B(\ImageBuffer[33][3] ), .C(
        \ImageBuffer[34][3] ), .D(\ImageBuffer[35][3] ), .S0(n3498), .S1(n3749), .Y(n3641) );
  MX4X1 U6551 ( .A(\ImageBuffer[0][6] ), .B(\ImageBuffer[1][6] ), .C(
        \ImageBuffer[2][6] ), .D(\ImageBuffer[3][6] ), .S0(n3488), .S1(n4130), 
        .Y(n3711) );
  MX4X1 U6552 ( .A(\ImageBuffer[32][6] ), .B(\ImageBuffer[33][6] ), .C(
        \ImageBuffer[34][6] ), .D(\ImageBuffer[35][6] ), .S0(n4116), .S1(n3749), .Y(n3701) );
  MX4X1 U6553 ( .A(\ImageBuffer[16][6] ), .B(\ImageBuffer[17][6] ), .C(
        \ImageBuffer[18][6] ), .D(\ImageBuffer[19][6] ), .S0(n4115), .S1(n4128), .Y(n3706) );
  MX4X1 U6554 ( .A(\ImageBuffer[48][6] ), .B(\ImageBuffer[49][6] ), .C(
        \ImageBuffer[50][6] ), .D(\ImageBuffer[51][6] ), .S0(n3743), .S1(n3753), .Y(n3696) );
  MX4X1 U6555 ( .A(\ImageBuffer[0][5] ), .B(\ImageBuffer[1][5] ), .C(
        \ImageBuffer[2][5] ), .D(\ImageBuffer[3][5] ), .S0(n4117), .S1(n3752), 
        .Y(n4066) );
  MX4X1 U6556 ( .A(\ImageBuffer[0][6] ), .B(\ImageBuffer[1][6] ), .C(
        \ImageBuffer[2][6] ), .D(\ImageBuffer[3][6] ), .S0(n4118), .S1(N2494), 
        .Y(n4086) );
  MX4X1 U6557 ( .A(\ImageBuffer[16][3] ), .B(\ImageBuffer[17][3] ), .C(
        \ImageBuffer[18][3] ), .D(\ImageBuffer[19][3] ), .S0(n3489), .S1(n3921), .Y(n3833) );
  MX4X1 U6558 ( .A(\ImageBuffer[48][3] ), .B(\ImageBuffer[49][3] ), .C(
        \ImageBuffer[50][3] ), .D(\ImageBuffer[51][3] ), .S0(n3489), .S1(n3480), .Y(n3823) );
  MX4X1 U6559 ( .A(\ImageBuffer[32][3] ), .B(\ImageBuffer[33][3] ), .C(
        \ImageBuffer[34][3] ), .D(\ImageBuffer[35][3] ), .S0(n3489), .S1(n3929), .Y(n3828) );
  MX4X1 U6560 ( .A(\ImageBuffer[32][4] ), .B(\ImageBuffer[33][4] ), .C(
        \ImageBuffer[34][4] ), .D(\ImageBuffer[35][4] ), .S0(n3742), .S1(n4129), .Y(n3661) );
  MX4X1 U6561 ( .A(\ImageBuffer[0][4] ), .B(\ImageBuffer[1][4] ), .C(
        \ImageBuffer[2][4] ), .D(\ImageBuffer[3][4] ), .S0(n4116), .S1(n3756), 
        .Y(n3671) );
  MX4X1 U6562 ( .A(\ImageBuffer[16][4] ), .B(\ImageBuffer[17][4] ), .C(
        \ImageBuffer[18][4] ), .D(\ImageBuffer[19][4] ), .S0(n3486), .S1(n3922), .Y(n3853) );
  MX4X1 U6563 ( .A(\ImageBuffer[48][4] ), .B(\ImageBuffer[49][4] ), .C(
        \ImageBuffer[50][4] ), .D(\ImageBuffer[51][4] ), .S0(n3486), .S1(n3932), .Y(n3843) );
  MX4X1 U6564 ( .A(\ImageBuffer[32][4] ), .B(\ImageBuffer[33][4] ), .C(
        \ImageBuffer[34][4] ), .D(\ImageBuffer[35][4] ), .S0(n3486), .S1(n3920), .Y(n3848) );
  MX4X1 U6565 ( .A(\ImageBuffer[0][4] ), .B(\ImageBuffer[1][4] ), .C(
        \ImageBuffer[2][4] ), .D(\ImageBuffer[3][4] ), .S0(n3941), .S1(n3929), 
        .Y(n3858) );
  MX4X1 U6566 ( .A(\ImageBuffer[48][2] ), .B(\ImageBuffer[49][2] ), .C(
        \ImageBuffer[50][2] ), .D(\ImageBuffer[51][2] ), .S0(n4300), .S1(n4312), .Y(n4180) );
  MX4X1 U6567 ( .A(\ImageBuffer[0][2] ), .B(\ImageBuffer[1][2] ), .C(
        \ImageBuffer[2][2] ), .D(\ImageBuffer[3][2] ), .S0(n3938), .S1(n4309), 
        .Y(n4195) );
  MX4X1 U6568 ( .A(\ImageBuffer[32][2] ), .B(\ImageBuffer[33][2] ), .C(
        \ImageBuffer[34][2] ), .D(\ImageBuffer[35][2] ), .S0(n3938), .S1(n4305), .Y(n4185) );
  MX4X1 U6569 ( .A(\ImageBuffer[32][6] ), .B(\ImageBuffer[33][6] ), .C(
        \ImageBuffer[34][6] ), .D(\ImageBuffer[35][6] ), .S0(n3939), .S1(n5123), .Y(n3888) );
  MX4X1 U6570 ( .A(\ImageBuffer[0][4] ), .B(\ImageBuffer[1][4] ), .C(
        \ImageBuffer[2][4] ), .D(\ImageBuffer[3][4] ), .S0(n3939), .S1(n4303), 
        .Y(n4235) );
  MX4X1 U6571 ( .A(\ImageBuffer[32][4] ), .B(\ImageBuffer[33][4] ), .C(
        \ImageBuffer[34][4] ), .D(\ImageBuffer[35][4] ), .S0(n3939), .S1(n4303), .Y(n4225) );
  MX4X1 U6572 ( .A(\ImageBuffer[16][4] ), .B(\ImageBuffer[17][4] ), .C(
        \ImageBuffer[18][4] ), .D(\ImageBuffer[19][4] ), .S0(n3941), .S1(n4309), .Y(n4230) );
  MX4X1 U6573 ( .A(\ImageBuffer[48][4] ), .B(\ImageBuffer[49][4] ), .C(
        \ImageBuffer[50][4] ), .D(\ImageBuffer[51][4] ), .S0(n4300), .S1(n5113), .Y(n4220) );
  MX4X1 U6574 ( .A(\ImageBuffer[0][6] ), .B(\ImageBuffer[1][6] ), .C(
        \ImageBuffer[2][6] ), .D(\ImageBuffer[3][6] ), .S0(n4297), .S1(n4307), 
        .Y(n4275) );
  MX4X1 U6575 ( .A(\ImageBuffer[32][6] ), .B(\ImageBuffer[33][6] ), .C(
        \ImageBuffer[34][6] ), .D(\ImageBuffer[35][6] ), .S0(n4297), .S1(n4303), .Y(n4265) );
  MX4X1 U6576 ( .A(\ImageBuffer[16][0] ), .B(\ImageBuffer[17][0] ), .C(
        \ImageBuffer[18][0] ), .D(\ImageBuffer[19][0] ), .S0(n3939), .S1(n4305), .Y(n4150) );
  MX4X1 U6577 ( .A(\ImageBuffer[48][0] ), .B(\ImageBuffer[49][0] ), .C(
        \ImageBuffer[50][0] ), .D(\ImageBuffer[51][0] ), .S0(n3939), .S1(n4307), .Y(n4140) );
  MX4X1 U6578 ( .A(\ImageBuffer[0][0] ), .B(\ImageBuffer[1][0] ), .C(
        \ImageBuffer[2][0] ), .D(\ImageBuffer[3][0] ), .S0(n3939), .S1(n4308), 
        .Y(n4155) );
  MX4X1 U6579 ( .A(\ImageBuffer[32][0] ), .B(\ImageBuffer[33][0] ), .C(
        \ImageBuffer[34][0] ), .D(\ImageBuffer[35][0] ), .S0(n3939), .S1(n5113), .Y(n4145) );
  MX4X1 U6580 ( .A(\ImageBuffer[0][0] ), .B(\ImageBuffer[1][0] ), .C(
        \ImageBuffer[2][0] ), .D(\ImageBuffer[3][0] ), .S0(n3512), .S1(n3472), 
        .Y(n4337) );
  MX4X1 U6581 ( .A(\ImageBuffer[32][0] ), .B(\ImageBuffer[33][0] ), .C(
        \ImageBuffer[34][0] ), .D(\ImageBuffer[35][0] ), .S0(n3514), .S1(n3473), .Y(n4327) );
  MX4X1 U6582 ( .A(\ImageBuffer[16][1] ), .B(\ImageBuffer[17][1] ), .C(
        \ImageBuffer[18][1] ), .D(\ImageBuffer[19][1] ), .S0(n3347), .S1(n3485), .Y(n4512) );
  MX4X1 U6583 ( .A(\ImageBuffer[32][1] ), .B(\ImageBuffer[33][1] ), .C(
        \ImageBuffer[34][1] ), .D(\ImageBuffer[35][1] ), .S0(n3343), .S1(n3485), .Y(n4507) );
  MX4X1 U6584 ( .A(\ImageBuffer[0][1] ), .B(\ImageBuffer[1][1] ), .C(
        \ImageBuffer[2][1] ), .D(\ImageBuffer[3][1] ), .S0(n3506), .S1(n3482), 
        .Y(n4517) );
  MX4X1 U6585 ( .A(\ImageBuffer[16][3] ), .B(\ImageBuffer[17][3] ), .C(
        \ImageBuffer[18][3] ), .D(\ImageBuffer[19][3] ), .S0(n3512), .S1(n3473), .Y(n4392) );
  MX4X1 U6586 ( .A(\ImageBuffer[32][3] ), .B(\ImageBuffer[33][3] ), .C(
        \ImageBuffer[34][3] ), .D(\ImageBuffer[35][3] ), .S0(n3511), .S1(n3474), .Y(n4387) );
  MX4X1 U6587 ( .A(\ImageBuffer[48][4] ), .B(\ImageBuffer[49][4] ), .C(
        \ImageBuffer[50][4] ), .D(\ImageBuffer[51][4] ), .S0(n3511), .S1(n3473), .Y(n4402) );
  MX4X1 U6588 ( .A(\ImageBuffer[32][4] ), .B(\ImageBuffer[33][4] ), .C(
        \ImageBuffer[34][4] ), .D(\ImageBuffer[35][4] ), .S0(n3515), .S1(n3472), .Y(n4407) );
  MX4X1 U6589 ( .A(\ImageBuffer[0][4] ), .B(\ImageBuffer[1][4] ), .C(
        \ImageBuffer[2][4] ), .D(\ImageBuffer[3][4] ), .S0(n3517), .S1(n3474), 
        .Y(n4417) );
  MX4X1 U6590 ( .A(\ImageBuffer[48][5] ), .B(\ImageBuffer[49][5] ), .C(
        \ImageBuffer[50][5] ), .D(\ImageBuffer[51][5] ), .S0(n3512), .S1(n3472), .Y(n4422) );
  MX4X1 U6591 ( .A(\ImageBuffer[32][5] ), .B(\ImageBuffer[33][5] ), .C(
        \ImageBuffer[34][5] ), .D(\ImageBuffer[35][5] ), .S0(n3518), .S1(n3472), .Y(n4427) );
  MX4X1 U6592 ( .A(\ImageBuffer[0][5] ), .B(\ImageBuffer[1][5] ), .C(
        \ImageBuffer[2][5] ), .D(\ImageBuffer[3][5] ), .S0(n3519), .S1(n3473), 
        .Y(n4437) );
  MX4X1 U6593 ( .A(\ImageBuffer[48][6] ), .B(\ImageBuffer[49][6] ), .C(
        \ImageBuffer[50][6] ), .D(\ImageBuffer[51][6] ), .S0(n3516), .S1(n3471), .Y(n4442) );
  MX4X1 U6594 ( .A(\ImageBuffer[32][6] ), .B(\ImageBuffer[33][6] ), .C(
        \ImageBuffer[34][6] ), .D(\ImageBuffer[35][6] ), .S0(n3512), .S1(n3473), .Y(n4447) );
  MX4X1 U6595 ( .A(\ImageBuffer[0][6] ), .B(\ImageBuffer[1][6] ), .C(
        \ImageBuffer[2][6] ), .D(\ImageBuffer[3][6] ), .S0(n3513), .S1(n3472), 
        .Y(n4457) );
  MX4X1 U6596 ( .A(\ImageBuffer[48][6] ), .B(\ImageBuffer[49][6] ), .C(
        \ImageBuffer[50][6] ), .D(\ImageBuffer[51][6] ), .S0(n3506), .S1(n3482), .Y(n4602) );
  MX4X1 U6597 ( .A(\ImageBuffer[32][6] ), .B(\ImageBuffer[33][6] ), .C(
        \ImageBuffer[34][6] ), .D(\ImageBuffer[35][6] ), .S0(n3506), .S1(n3482), .Y(n4607) );
  MX4X1 U6598 ( .A(\ImageBuffer[0][6] ), .B(\ImageBuffer[1][6] ), .C(
        \ImageBuffer[2][6] ), .D(\ImageBuffer[3][6] ), .S0(n3347), .S1(n3484), 
        .Y(n4617) );
  MX4X1 U6599 ( .A(\ImageBuffer[48][7] ), .B(\ImageBuffer[49][7] ), .C(
        \ImageBuffer[50][7] ), .D(\ImageBuffer[51][7] ), .S0(n3519), .S1(n3473), .Y(n4462) );
  MX4X1 U6600 ( .A(\ImageBuffer[32][7] ), .B(\ImageBuffer[33][7] ), .C(
        \ImageBuffer[34][7] ), .D(\ImageBuffer[35][7] ), .S0(n3511), .S1(n3474), .Y(n4467) );
  MX4X1 U6601 ( .A(\ImageBuffer[0][7] ), .B(\ImageBuffer[1][7] ), .C(
        \ImageBuffer[2][7] ), .D(\ImageBuffer[3][7] ), .S0(n3513), .S1(n3472), 
        .Y(n4477) );
  MX4X1 U6602 ( .A(\ImageBuffer[48][7] ), .B(\ImageBuffer[49][7] ), .C(
        \ImageBuffer[50][7] ), .D(\ImageBuffer[51][7] ), .S0(n3342), .S1(n3485), .Y(n4622) );
  MX4X1 U6603 ( .A(\ImageBuffer[32][7] ), .B(\ImageBuffer[33][7] ), .C(
        \ImageBuffer[34][7] ), .D(\ImageBuffer[35][7] ), .S0(n3346), .S1(n3484), .Y(n4627) );
  MX4X1 U6604 ( .A(\ImageBuffer[0][7] ), .B(\ImageBuffer[1][7] ), .C(
        \ImageBuffer[2][7] ), .D(\ImageBuffer[3][7] ), .S0(n3506), .S1(n3483), 
        .Y(n4637) );
  MX4X1 U6605 ( .A(\ImageBuffer[32][4] ), .B(\ImageBuffer[33][4] ), .C(
        \ImageBuffer[34][4] ), .D(\ImageBuffer[35][4] ), .S0(n4119), .S1(n3749), .Y(n4036) );
  MX4X1 U6606 ( .A(\ImageBuffer[0][4] ), .B(\ImageBuffer[1][4] ), .C(
        \ImageBuffer[2][4] ), .D(\ImageBuffer[3][4] ), .S0(n4116), .S1(n4123), 
        .Y(n4046) );
  MX4X1 U6607 ( .A(\ImageBuffer[24][0] ), .B(\ImageBuffer[25][0] ), .C(
        \ImageBuffer[26][0] ), .D(\ImageBuffer[27][0] ), .S0(n3742), .S1(n3750), .Y(n3584) );
  MX4X1 U6608 ( .A(\ImageBuffer[28][0] ), .B(\ImageBuffer[29][0] ), .C(
        \ImageBuffer[30][0] ), .D(\ImageBuffer[31][0] ), .S0(n3742), .S1(n4127), .Y(n3583) );
  MX4X1 U6609 ( .A(\ImageBuffer[20][0] ), .B(\ImageBuffer[21][0] ), .C(
        \ImageBuffer[22][0] ), .D(\ImageBuffer[23][0] ), .S0(n3742), .S1(n4134), .Y(n3585) );
  MX4X1 U6610 ( .A(\ImageBuffer[24][0] ), .B(\ImageBuffer[25][0] ), .C(
        \ImageBuffer[26][0] ), .D(\ImageBuffer[27][0] ), .S0(n3938), .S1(n3341), .Y(n3771) );
  MX4X1 U6611 ( .A(\ImageBuffer[28][0] ), .B(\ImageBuffer[29][0] ), .C(
        \ImageBuffer[30][0] ), .D(\ImageBuffer[31][0] ), .S0(n3938), .S1(n3927), .Y(n3770) );
  MX4X1 U6612 ( .A(\ImageBuffer[20][0] ), .B(\ImageBuffer[21][0] ), .C(
        \ImageBuffer[22][0] ), .D(\ImageBuffer[23][0] ), .S0(n3938), .S1(n3927), .Y(n3772) );
  MX4X1 U6613 ( .A(\ImageBuffer[24][0] ), .B(\ImageBuffer[25][0] ), .C(
        \ImageBuffer[26][0] ), .D(\ImageBuffer[27][0] ), .S0(n3506), .S1(n3484), .Y(n4490) );
  MX4X1 U6614 ( .A(\ImageBuffer[28][0] ), .B(\ImageBuffer[29][0] ), .C(
        \ImageBuffer[30][0] ), .D(\ImageBuffer[31][0] ), .S0(n3343), .S1(n3483), .Y(n4489) );
  MX4X1 U6615 ( .A(\ImageBuffer[20][0] ), .B(\ImageBuffer[21][0] ), .C(
        \ImageBuffer[22][0] ), .D(\ImageBuffer[23][0] ), .S0(n3347), .S1(n3482), .Y(n4491) );
  MX4X1 U6616 ( .A(\ImageBuffer[16][2] ), .B(\ImageBuffer[17][2] ), .C(
        \ImageBuffer[18][2] ), .D(\ImageBuffer[19][2] ), .S0(n3939), .S1(n3932), .Y(n3813) );
  MX4X1 U6617 ( .A(\ImageBuffer[24][2] ), .B(\ImageBuffer[25][2] ), .C(
        \ImageBuffer[26][2] ), .D(\ImageBuffer[27][2] ), .S0(n3939), .S1(n3340), .Y(n3811) );
  MX4X1 U6618 ( .A(\ImageBuffer[28][2] ), .B(\ImageBuffer[29][2] ), .C(
        \ImageBuffer[30][2] ), .D(\ImageBuffer[31][2] ), .S0(n3939), .S1(n3930), .Y(n3810) );
  MX4X1 U6619 ( .A(n3626), .B(n3624), .C(n3625), .D(n3623), .S0(n3734), .S1(
        n3758), .Y(n3627) );
  MX4X1 U6620 ( .A(\ImageBuffer[16][2] ), .B(\ImageBuffer[17][2] ), .C(
        \ImageBuffer[18][2] ), .D(\ImageBuffer[19][2] ), .S0(n3741), .S1(n4126), .Y(n3626) );
  MX4X1 U6621 ( .A(\ImageBuffer[24][2] ), .B(\ImageBuffer[25][2] ), .C(
        \ImageBuffer[26][2] ), .D(\ImageBuffer[27][2] ), .S0(n3741), .S1(n3753), .Y(n3624) );
  MX4X1 U6622 ( .A(\ImageBuffer[28][2] ), .B(\ImageBuffer[29][2] ), .C(
        \ImageBuffer[30][2] ), .D(\ImageBuffer[31][2] ), .S0(n3741), .S1(n3751), .Y(n3623) );
  MX4X1 U6623 ( .A(\ImageBuffer[16][3] ), .B(\ImageBuffer[17][3] ), .C(
        \ImageBuffer[18][3] ), .D(\ImageBuffer[19][3] ), .S0(n3498), .S1(n3753), .Y(n3646) );
  MX4X1 U6624 ( .A(\ImageBuffer[24][3] ), .B(\ImageBuffer[25][3] ), .C(
        \ImageBuffer[26][3] ), .D(\ImageBuffer[27][3] ), .S0(n3498), .S1(n4123), .Y(n3644) );
  MX4X1 U6625 ( .A(\ImageBuffer[28][3] ), .B(\ImageBuffer[29][3] ), .C(
        \ImageBuffer[30][3] ), .D(\ImageBuffer[31][3] ), .S0(n3498), .S1(n3754), .Y(n3643) );
  MX4X1 U6626 ( .A(n4061), .B(n4059), .C(n4060), .D(n4058), .S0(n4109), .S1(
        n4136), .Y(n4062) );
  MX4X1 U6627 ( .A(\ImageBuffer[16][5] ), .B(\ImageBuffer[17][5] ), .C(
        \ImageBuffer[18][5] ), .D(\ImageBuffer[19][5] ), .S0(n4117), .S1(n3749), .Y(n4061) );
  MX4X1 U6628 ( .A(\ImageBuffer[24][5] ), .B(\ImageBuffer[25][5] ), .C(
        \ImageBuffer[26][5] ), .D(\ImageBuffer[27][5] ), .S0(n4117), .S1(n3747), .Y(n4059) );
  MX4X1 U6629 ( .A(n4081), .B(n4079), .C(n4080), .D(n4078), .S0(n4109), .S1(
        n4136), .Y(n4082) );
  MX4X1 U6630 ( .A(\ImageBuffer[16][6] ), .B(\ImageBuffer[17][6] ), .C(
        \ImageBuffer[18][6] ), .D(\ImageBuffer[19][6] ), .S0(n4118), .S1(n4123), .Y(n4081) );
  MX4X1 U6631 ( .A(\ImageBuffer[24][6] ), .B(\ImageBuffer[25][6] ), .C(
        \ImageBuffer[26][6] ), .D(\ImageBuffer[27][6] ), .S0(n4118), .S1(n4128), .Y(n4079) );
  MX4X1 U6632 ( .A(\ImageBuffer[24][3] ), .B(\ImageBuffer[25][3] ), .C(
        \ImageBuffer[26][3] ), .D(\ImageBuffer[27][3] ), .S0(n4116), .S1(n4129), .Y(n4019) );
  MX4X1 U6633 ( .A(\ImageBuffer[28][3] ), .B(\ImageBuffer[29][3] ), .C(
        \ImageBuffer[30][3] ), .D(\ImageBuffer[31][3] ), .S0(n4116), .S1(n3754), .Y(n4018) );
  MX4X1 U6634 ( .A(n3666), .B(n3664), .C(n3665), .D(n3663), .S0(n3734), .S1(
        n3758), .Y(n3667) );
  MX4X1 U6635 ( .A(\ImageBuffer[16][4] ), .B(\ImageBuffer[17][4] ), .C(
        \ImageBuffer[18][4] ), .D(\ImageBuffer[19][4] ), .S0(n3742), .S1(n4128), .Y(n3666) );
  MX4X1 U6636 ( .A(n4270), .B(n4268), .C(n4269), .D(n4267), .S0(n5108), .S1(
        n3487), .Y(n4271) );
  MX4X1 U6637 ( .A(\ImageBuffer[16][6] ), .B(\ImageBuffer[17][6] ), .C(
        \ImageBuffer[18][6] ), .D(\ImageBuffer[19][6] ), .S0(n3935), .S1(n4315), .Y(n4270) );
  MX4X1 U6638 ( .A(\ImageBuffer[24][6] ), .B(\ImageBuffer[25][6] ), .C(
        \ImageBuffer[26][6] ), .D(\ImageBuffer[27][6] ), .S0(n3935), .S1(n4311), .Y(n4268) );
  MX4X1 U6639 ( .A(\ImageBuffer[28][6] ), .B(\ImageBuffer[29][6] ), .C(
        \ImageBuffer[30][6] ), .D(\ImageBuffer[31][6] ), .S0(n4297), .S1(n4314), .Y(n4267) );
  MX4X1 U6640 ( .A(\ImageBuffer[16][7] ), .B(\ImageBuffer[17][7] ), .C(
        \ImageBuffer[18][7] ), .D(\ImageBuffer[19][7] ), .S0(n3939), .S1(n4317), .Y(n4290) );
  MX4X1 U6641 ( .A(\ImageBuffer[24][7] ), .B(\ImageBuffer[25][7] ), .C(
        \ImageBuffer[26][7] ), .D(\ImageBuffer[27][7] ), .S0(n3939), .S1(n4309), .Y(n4288) );
  MX4X1 U6642 ( .A(\ImageBuffer[28][7] ), .B(\ImageBuffer[29][7] ), .C(
        \ImageBuffer[30][7] ), .D(\ImageBuffer[31][7] ), .S0(n3939), .S1(n4313), .Y(n4287) );
  MX4X1 U6643 ( .A(\ImageBuffer[16][1] ), .B(\ImageBuffer[17][1] ), .C(
        \ImageBuffer[18][1] ), .D(\ImageBuffer[19][1] ), .S0(n3522), .S1(n3473), .Y(n4352) );
  MX4X1 U6644 ( .A(\ImageBuffer[24][1] ), .B(\ImageBuffer[25][1] ), .C(
        \ImageBuffer[26][1] ), .D(\ImageBuffer[27][1] ), .S0(n3521), .S1(n3472), .Y(n4350) );
  MX4X1 U6645 ( .A(n4552), .B(n4550), .C(n4551), .D(n4549), .S0(n3496), .S1(
        n4639), .Y(n4553) );
  MX4X1 U6646 ( .A(\ImageBuffer[16][3] ), .B(\ImageBuffer[17][3] ), .C(
        \ImageBuffer[18][3] ), .D(\ImageBuffer[19][3] ), .S0(n3343), .S1(n3483), .Y(n4552) );
  MX4X1 U6647 ( .A(\ImageBuffer[24][3] ), .B(\ImageBuffer[25][3] ), .C(
        \ImageBuffer[26][3] ), .D(\ImageBuffer[27][3] ), .S0(n3347), .S1(n3484), .Y(n4550) );
  MX4X1 U6648 ( .A(\ImageBuffer[28][3] ), .B(\ImageBuffer[29][3] ), .C(
        \ImageBuffer[30][3] ), .D(\ImageBuffer[31][3] ), .S0(n3347), .S1(n3483), .Y(n4549) );
  MX4X1 U6649 ( .A(n4412), .B(n4410), .C(n4411), .D(n4409), .S0(n3503), .S1(
        n3495), .Y(n4413) );
  MX4X1 U6650 ( .A(\ImageBuffer[16][4] ), .B(\ImageBuffer[17][4] ), .C(
        \ImageBuffer[18][4] ), .D(\ImageBuffer[19][4] ), .S0(n3513), .S1(n3471), .Y(n4412) );
  MX4X1 U6651 ( .A(\ImageBuffer[24][4] ), .B(\ImageBuffer[25][4] ), .C(
        \ImageBuffer[26][4] ), .D(\ImageBuffer[27][4] ), .S0(n3511), .S1(n3473), .Y(n4410) );
  MX4X1 U6652 ( .A(\ImageBuffer[28][4] ), .B(\ImageBuffer[29][4] ), .C(
        \ImageBuffer[30][4] ), .D(\ImageBuffer[31][4] ), .S0(n3521), .S1(n3474), .Y(n4409) );
  MX4X1 U6653 ( .A(n4432), .B(n4430), .C(n4431), .D(n4429), .S0(n3503), .S1(
        n3495), .Y(n4433) );
  MX4X1 U6654 ( .A(\ImageBuffer[16][5] ), .B(\ImageBuffer[17][5] ), .C(
        \ImageBuffer[18][5] ), .D(\ImageBuffer[19][5] ), .S0(n3514), .S1(n3474), .Y(n4432) );
  MX4X1 U6655 ( .A(\ImageBuffer[24][5] ), .B(\ImageBuffer[25][5] ), .C(
        \ImageBuffer[26][5] ), .D(\ImageBuffer[27][5] ), .S0(n3513), .S1(n3471), .Y(n4430) );
  MX4X1 U6656 ( .A(\ImageBuffer[28][5] ), .B(\ImageBuffer[29][5] ), .C(
        \ImageBuffer[30][5] ), .D(\ImageBuffer[31][5] ), .S0(n3511), .S1(n3474), .Y(n4429) );
  MX4X1 U6657 ( .A(n4472), .B(n4470), .C(n4471), .D(n4469), .S0(n3503), .S1(
        n3495), .Y(n4473) );
  MX4X1 U6658 ( .A(\ImageBuffer[16][7] ), .B(\ImageBuffer[17][7] ), .C(
        \ImageBuffer[18][7] ), .D(\ImageBuffer[19][7] ), .S0(n3513), .S1(n3473), .Y(n4472) );
  MX4X1 U6659 ( .A(\ImageBuffer[24][7] ), .B(\ImageBuffer[25][7] ), .C(
        \ImageBuffer[26][7] ), .D(\ImageBuffer[27][7] ), .S0(n3512), .S1(n3471), .Y(n4470) );
  MX4X1 U6660 ( .A(\ImageBuffer[28][7] ), .B(\ImageBuffer[29][7] ), .C(
        \ImageBuffer[30][7] ), .D(\ImageBuffer[31][7] ), .S0(n3511), .S1(n3473), .Y(n4469) );
  MX4X1 U6661 ( .A(\ImageBuffer[16][4] ), .B(\ImageBuffer[17][4] ), .C(
        \ImageBuffer[18][4] ), .D(\ImageBuffer[19][4] ), .S0(n4119), .S1(n4122), .Y(n4041) );
  MX4X1 U6662 ( .A(\ImageBuffer[24][4] ), .B(\ImageBuffer[25][4] ), .C(
        \ImageBuffer[26][4] ), .D(\ImageBuffer[27][4] ), .S0(n4119), .S1(n4130), .Y(n4039) );
  MX4X1 U6663 ( .A(\ImageBuffer[28][4] ), .B(\ImageBuffer[29][4] ), .C(
        \ImageBuffer[30][4] ), .D(\ImageBuffer[31][4] ), .S0(n4119), .S1(n4128), .Y(n4038) );
  MX4X1 U6664 ( .A(n3591), .B(n3589), .C(n3590), .D(n3588), .S0(n3733), .S1(
        n3758), .Y(n3592) );
  MX4X1 U6665 ( .A(\ImageBuffer[0][0] ), .B(\ImageBuffer[1][0] ), .C(
        \ImageBuffer[2][0] ), .D(\ImageBuffer[3][0] ), .S0(n3740), .S1(n3749), 
        .Y(n3591) );
  MX4X1 U6666 ( .A(\ImageBuffer[8][0] ), .B(\ImageBuffer[9][0] ), .C(
        \ImageBuffer[10][0] ), .D(\ImageBuffer[11][0] ), .S0(n3740), .S1(n4130), .Y(n3589) );
  MX4X1 U6667 ( .A(\ImageBuffer[12][0] ), .B(\ImageBuffer[13][0] ), .C(
        \ImageBuffer[14][0] ), .D(\ImageBuffer[15][0] ), .S0(n3740), .S1(n4130), .Y(n3588) );
  MX4X1 U6668 ( .A(\ImageBuffer[0][0] ), .B(\ImageBuffer[1][0] ), .C(
        \ImageBuffer[2][0] ), .D(\ImageBuffer[3][0] ), .S0(n3939), .S1(n3924), 
        .Y(n3778) );
  MX4X1 U6669 ( .A(\ImageBuffer[8][0] ), .B(\ImageBuffer[9][0] ), .C(
        \ImageBuffer[10][0] ), .D(\ImageBuffer[11][0] ), .S0(n3939), .S1(n5123), .Y(n3776) );
  MX4X1 U6670 ( .A(\ImageBuffer[12][0] ), .B(\ImageBuffer[13][0] ), .C(
        \ImageBuffer[14][0] ), .D(\ImageBuffer[15][0] ), .S0(n3939), .S1(n3921), .Y(n3775) );
  MX4X1 U6671 ( .A(n4497), .B(n4495), .C(n4496), .D(n4494), .S0(n3496), .S1(
        n4641), .Y(n4498) );
  MX4X1 U6672 ( .A(\ImageBuffer[0][0] ), .B(\ImageBuffer[1][0] ), .C(
        \ImageBuffer[2][0] ), .D(\ImageBuffer[3][0] ), .S0(n3343), .S1(n3485), 
        .Y(n4497) );
  MX4X1 U6673 ( .A(\ImageBuffer[8][0] ), .B(\ImageBuffer[9][0] ), .C(
        \ImageBuffer[10][0] ), .D(\ImageBuffer[11][0] ), .S0(n3347), .S1(n3483), .Y(n4495) );
  MX4X1 U6674 ( .A(\ImageBuffer[12][0] ), .B(\ImageBuffer[13][0] ), .C(
        \ImageBuffer[14][0] ), .D(\ImageBuffer[15][0] ), .S0(n3343), .S1(n3485), .Y(n4494) );
  MX4X1 U6675 ( .A(\ImageBuffer[12][4] ), .B(\ImageBuffer[13][4] ), .C(
        \ImageBuffer[14][4] ), .D(\ImageBuffer[15][4] ), .S0(n3939), .S1(n4310), .Y(n4232) );
  MX4X1 U6676 ( .A(\ImageBuffer[4][4] ), .B(\ImageBuffer[5][4] ), .C(
        \ImageBuffer[6][4] ), .D(\ImageBuffer[7][4] ), .S0(n3939), .S1(n4313), 
        .Y(n4234) );
  MX4X1 U6677 ( .A(\ImageBuffer[8][4] ), .B(\ImageBuffer[9][4] ), .C(
        \ImageBuffer[10][4] ), .D(\ImageBuffer[11][4] ), .S0(n3939), .S1(n4313), .Y(n4233) );
  MX4X1 U6678 ( .A(n3711), .B(n3709), .C(n3710), .D(n3708), .S0(n3734), .S1(
        n3759), .Y(n3712) );
  MX4X1 U6679 ( .A(\ImageBuffer[12][6] ), .B(\ImageBuffer[13][6] ), .C(
        \ImageBuffer[14][6] ), .D(\ImageBuffer[15][6] ), .S0(n4115), .S1(n4129), .Y(n3708) );
  MX4X1 U6680 ( .A(\ImageBuffer[4][6] ), .B(\ImageBuffer[5][6] ), .C(
        \ImageBuffer[6][6] ), .D(\ImageBuffer[7][6] ), .S0(n4115), .S1(n4125), 
        .Y(n3710) );
  MX4X1 U6681 ( .A(\ImageBuffer[8][6] ), .B(\ImageBuffer[9][6] ), .C(
        \ImageBuffer[10][6] ), .D(\ImageBuffer[11][6] ), .S0(n4115), .S1(n3752), .Y(n3709) );
  MX4X1 U6682 ( .A(n4357), .B(n4355), .C(n4356), .D(n4354), .S0(n3503), .S1(
        n3495), .Y(n4358) );
  MX4X1 U6683 ( .A(\ImageBuffer[0][1] ), .B(\ImageBuffer[1][1] ), .C(
        \ImageBuffer[2][1] ), .D(\ImageBuffer[3][1] ), .S0(n3519), .S1(n3472), 
        .Y(n4357) );
  MX4X1 U6684 ( .A(\ImageBuffer[8][1] ), .B(\ImageBuffer[9][1] ), .C(
        \ImageBuffer[10][1] ), .D(\ImageBuffer[11][1] ), .S0(n3518), .S1(n3472), .Y(n4355) );
  MX4X1 U6685 ( .A(\ImageBuffer[12][1] ), .B(\ImageBuffer[13][1] ), .C(
        \ImageBuffer[14][1] ), .D(\ImageBuffer[15][1] ), .S0(n3514), .S1(n3471), .Y(n4354) );
  MX4X1 U6686 ( .A(n4557), .B(n4555), .C(n4556), .D(n4554), .S0(n3496), .S1(
        n4639), .Y(n4558) );
  MX4X1 U6687 ( .A(\ImageBuffer[8][3] ), .B(\ImageBuffer[9][3] ), .C(
        \ImageBuffer[10][3] ), .D(\ImageBuffer[11][3] ), .S0(n3347), .S1(n3485), .Y(n4555) );
  MX4X1 U6688 ( .A(\ImageBuffer[12][3] ), .B(\ImageBuffer[13][3] ), .C(
        \ImageBuffer[14][3] ), .D(\ImageBuffer[15][3] ), .S0(n3347), .S1(n3482), .Y(n4554) );
  MX4X1 U6689 ( .A(\ImageBuffer[28][3] ), .B(\ImageBuffer[29][3] ), .C(
        \ImageBuffer[30][3] ), .D(\ImageBuffer[31][3] ), .S0(n3521), .S1(n3474), .Y(n4389) );
  MX4X1 U6690 ( .A(\ImageBuffer[44][2] ), .B(\ImageBuffer[45][2] ), .C(
        \ImageBuffer[46][2] ), .D(\ImageBuffer[47][2] ), .S0(n4115), .S1(n3753), .Y(n3993) );
  MX4X1 U6691 ( .A(\ImageBuffer[12][2] ), .B(\ImageBuffer[13][2] ), .C(
        \ImageBuffer[14][2] ), .D(\ImageBuffer[15][2] ), .S0(n3735), .S1(n3748), .Y(n4003) );
  MX4X1 U6692 ( .A(\ImageBuffer[60][0] ), .B(\ImageBuffer[61][0] ), .C(
        \ImageBuffer[62][0] ), .D(\ImageBuffer[63][0] ), .S0(n4114), .S1(n4132), .Y(n3950) );
  MX4X1 U6693 ( .A(\ImageBuffer[44][0] ), .B(\ImageBuffer[45][0] ), .C(
        \ImageBuffer[46][0] ), .D(\ImageBuffer[47][0] ), .S0(n4114), .S1(n3747), .Y(n3954) );
  MX4X1 U6694 ( .A(\ImageBuffer[12][2] ), .B(\ImageBuffer[13][2] ), .C(
        \ImageBuffer[14][2] ), .D(\ImageBuffer[15][2] ), .S0(n3939), .S1(n3921), .Y(n3815) );
  MX4X1 U6695 ( .A(\ImageBuffer[60][0] ), .B(\ImageBuffer[61][0] ), .C(
        \ImageBuffer[62][0] ), .D(\ImageBuffer[63][0] ), .S0(n4117), .S1(n3755), .Y(n3573) );
  MX4X1 U6696 ( .A(\ImageBuffer[44][0] ), .B(\ImageBuffer[45][0] ), .C(
        \ImageBuffer[46][0] ), .D(\ImageBuffer[47][0] ), .S0(n4119), .S1(n4123), .Y(n3578) );
  MX4X1 U6697 ( .A(\ImageBuffer[28][0] ), .B(\ImageBuffer[29][0] ), .C(
        \ImageBuffer[30][0] ), .D(\ImageBuffer[31][0] ), .S0(n3517), .S1(n3471), .Y(n4329) );
  MX4X1 U6698 ( .A(\ImageBuffer[60][0] ), .B(\ImageBuffer[61][0] ), .C(
        \ImageBuffer[62][0] ), .D(\ImageBuffer[63][0] ), .S0(n3938), .S1(n3480), .Y(n3760) );
  MX4X1 U6699 ( .A(\ImageBuffer[44][0] ), .B(\ImageBuffer[45][0] ), .C(
        \ImageBuffer[46][0] ), .D(\ImageBuffer[47][0] ), .S0(n3938), .S1(n3925), .Y(n3765) );
  MX4X1 U6700 ( .A(\ImageBuffer[60][2] ), .B(\ImageBuffer[61][2] ), .C(
        \ImageBuffer[62][2] ), .D(\ImageBuffer[63][2] ), .S0(n3506), .S1(n3485), .Y(n4519) );
  MX4X1 U6701 ( .A(\ImageBuffer[44][2] ), .B(\ImageBuffer[45][2] ), .C(
        \ImageBuffer[46][2] ), .D(\ImageBuffer[47][2] ), .S0(n3347), .S1(n3485), .Y(n4524) );
  MX4X1 U6702 ( .A(\ImageBuffer[44][2] ), .B(\ImageBuffer[45][2] ), .C(
        \ImageBuffer[46][2] ), .D(\ImageBuffer[47][2] ), .S0(n3743), .S1(n4133), .Y(n3618) );
  MX4X1 U6703 ( .A(\ImageBuffer[12][2] ), .B(\ImageBuffer[13][2] ), .C(
        \ImageBuffer[14][2] ), .D(\ImageBuffer[15][2] ), .S0(n3741), .S1(n4129), .Y(n3628) );
  MX4X1 U6704 ( .A(\ImageBuffer[44][3] ), .B(\ImageBuffer[45][3] ), .C(
        \ImageBuffer[46][3] ), .D(\ImageBuffer[47][3] ), .S0(n3498), .S1(n4125), .Y(n3638) );
  MX4X1 U6705 ( .A(\ImageBuffer[12][3] ), .B(\ImageBuffer[13][3] ), .C(
        \ImageBuffer[14][3] ), .D(\ImageBuffer[15][3] ), .S0(n3498), .S1(n3755), .Y(n3648) );
  MX4X1 U6706 ( .A(\ImageBuffer[28][6] ), .B(\ImageBuffer[29][6] ), .C(
        \ImageBuffer[30][6] ), .D(\ImageBuffer[31][6] ), .S0(n4115), .S1(n4125), .Y(n3703) );
  MX4X1 U6707 ( .A(\ImageBuffer[60][6] ), .B(\ImageBuffer[61][6] ), .C(
        \ImageBuffer[62][6] ), .D(\ImageBuffer[63][6] ), .S0(n3743), .S1(n3752), .Y(n3693) );
  MX4X1 U6708 ( .A(\ImageBuffer[12][5] ), .B(\ImageBuffer[13][5] ), .C(
        \ImageBuffer[14][5] ), .D(\ImageBuffer[15][5] ), .S0(n4117), .S1(n4131), .Y(n4063) );
  MX4X1 U6709 ( .A(\ImageBuffer[12][3] ), .B(\ImageBuffer[13][3] ), .C(
        \ImageBuffer[14][3] ), .D(\ImageBuffer[15][3] ), .S0(n4116), .S1(n3749), .Y(n4023) );
  MX4X1 U6710 ( .A(\ImageBuffer[44][3] ), .B(\ImageBuffer[45][3] ), .C(
        \ImageBuffer[46][3] ), .D(\ImageBuffer[47][3] ), .S0(n3489), .S1(n3920), .Y(n3825) );
  MX4X1 U6711 ( .A(\ImageBuffer[44][4] ), .B(\ImageBuffer[45][4] ), .C(
        \ImageBuffer[46][4] ), .D(\ImageBuffer[47][4] ), .S0(n3742), .S1(n3750), .Y(n3658) );
  MX4X1 U6712 ( .A(\ImageBuffer[12][4] ), .B(\ImageBuffer[13][4] ), .C(
        \ImageBuffer[14][4] ), .D(\ImageBuffer[15][4] ), .S0(n3498), .S1(n4130), .Y(n3668) );
  MX4X1 U6713 ( .A(\ImageBuffer[44][4] ), .B(\ImageBuffer[45][4] ), .C(
        \ImageBuffer[46][4] ), .D(\ImageBuffer[47][4] ), .S0(n3486), .S1(n3921), .Y(n3845) );
  MX4X1 U6714 ( .A(\ImageBuffer[12][4] ), .B(\ImageBuffer[13][4] ), .C(
        \ImageBuffer[14][4] ), .D(\ImageBuffer[15][4] ), .S0(n4300), .S1(n3499), .Y(n3855) );
  MX4X1 U6715 ( .A(\ImageBuffer[60][2] ), .B(\ImageBuffer[61][2] ), .C(
        \ImageBuffer[62][2] ), .D(\ImageBuffer[63][2] ), .S0(n4300), .S1(n4306), .Y(n4177) );
  MX4X1 U6716 ( .A(\ImageBuffer[12][2] ), .B(\ImageBuffer[13][2] ), .C(
        \ImageBuffer[14][2] ), .D(\ImageBuffer[15][2] ), .S0(n3938), .S1(n4311), .Y(n4192) );
  MX4X1 U6717 ( .A(\ImageBuffer[44][2] ), .B(\ImageBuffer[45][2] ), .C(
        \ImageBuffer[46][2] ), .D(\ImageBuffer[47][2] ), .S0(n4300), .S1(n4309), .Y(n4182) );
  MX4X1 U6718 ( .A(\ImageBuffer[12][6] ), .B(\ImageBuffer[13][6] ), .C(
        \ImageBuffer[14][6] ), .D(\ImageBuffer[15][6] ), .S0(n3939), .S1(n3922), .Y(n3895) );
  MX4X1 U6719 ( .A(\ImageBuffer[44][4] ), .B(\ImageBuffer[45][4] ), .C(
        \ImageBuffer[46][4] ), .D(\ImageBuffer[47][4] ), .S0(n3935), .S1(n4315), .Y(n4222) );
  MX4X1 U6720 ( .A(\ImageBuffer[28][4] ), .B(\ImageBuffer[29][4] ), .C(
        \ImageBuffer[30][4] ), .D(\ImageBuffer[31][4] ), .S0(n3486), .S1(n4304), .Y(n4227) );
  MX4X1 U6721 ( .A(\ImageBuffer[60][4] ), .B(\ImageBuffer[61][4] ), .C(
        \ImageBuffer[62][4] ), .D(\ImageBuffer[63][4] ), .S0(n3940), .S1(n4308), .Y(n4217) );
  MX4X1 U6722 ( .A(\ImageBuffer[12][6] ), .B(\ImageBuffer[13][6] ), .C(
        \ImageBuffer[14][6] ), .D(\ImageBuffer[15][6] ), .S0(n3935), .S1(n4317), .Y(n4272) );
  MX4X1 U6723 ( .A(\ImageBuffer[60][0] ), .B(\ImageBuffer[61][0] ), .C(
        \ImageBuffer[62][0] ), .D(\ImageBuffer[63][0] ), .S0(n3938), .S1(n4304), .Y(n4137) );
  MX4X1 U6724 ( .A(\ImageBuffer[12][0] ), .B(\ImageBuffer[13][0] ), .C(
        \ImageBuffer[14][0] ), .D(\ImageBuffer[15][0] ), .S0(n3939), .S1(n4305), .Y(n4152) );
  MX4X1 U6725 ( .A(\ImageBuffer[44][0] ), .B(\ImageBuffer[45][0] ), .C(
        \ImageBuffer[46][0] ), .D(\ImageBuffer[47][0] ), .S0(n3938), .S1(n4313), .Y(n4142) );
  MX4X1 U6726 ( .A(\ImageBuffer[12][0] ), .B(\ImageBuffer[13][0] ), .C(
        \ImageBuffer[14][0] ), .D(\ImageBuffer[15][0] ), .S0(n3522), .S1(n3473), .Y(n4334) );
  MX4X1 U6727 ( .A(\ImageBuffer[44][0] ), .B(\ImageBuffer[45][0] ), .C(
        \ImageBuffer[46][0] ), .D(\ImageBuffer[47][0] ), .S0(n3514), .S1(n3473), .Y(n4324) );
  MX4X1 U6728 ( .A(\ImageBuffer[28][1] ), .B(\ImageBuffer[29][1] ), .C(
        \ImageBuffer[30][1] ), .D(\ImageBuffer[31][1] ), .S0(n3343), .S1(n3485), .Y(n4509) );
  MX4X1 U6729 ( .A(\ImageBuffer[44][1] ), .B(\ImageBuffer[45][1] ), .C(
        \ImageBuffer[46][1] ), .D(\ImageBuffer[47][1] ), .S0(n3343), .S1(n3483), .Y(n4504) );
  MX4X1 U6730 ( .A(\ImageBuffer[12][1] ), .B(\ImageBuffer[13][1] ), .C(
        \ImageBuffer[14][1] ), .D(\ImageBuffer[15][1] ), .S0(n3347), .S1(n3484), .Y(n4514) );
  MX4X1 U6731 ( .A(\ImageBuffer[44][3] ), .B(\ImageBuffer[45][3] ), .C(
        \ImageBuffer[46][3] ), .D(\ImageBuffer[47][3] ), .S0(n3511), .S1(n3473), .Y(n4384) );
  MX4X1 U6732 ( .A(\ImageBuffer[12][3] ), .B(\ImageBuffer[13][3] ), .C(
        \ImageBuffer[14][3] ), .D(\ImageBuffer[15][3] ), .S0(n3513), .S1(n3473), .Y(n4394) );
  MX4X1 U6733 ( .A(\ImageBuffer[60][4] ), .B(\ImageBuffer[61][4] ), .C(
        \ImageBuffer[62][4] ), .D(\ImageBuffer[63][4] ), .S0(n3512), .S1(n3471), .Y(n4399) );
  MX4X1 U6734 ( .A(\ImageBuffer[44][4] ), .B(\ImageBuffer[45][4] ), .C(
        \ImageBuffer[46][4] ), .D(\ImageBuffer[47][4] ), .S0(n3518), .S1(n3471), .Y(n4404) );
  MX4X1 U6735 ( .A(\ImageBuffer[12][4] ), .B(\ImageBuffer[13][4] ), .C(
        \ImageBuffer[14][4] ), .D(\ImageBuffer[15][4] ), .S0(n3521), .S1(n3471), .Y(n4414) );
  MX4X1 U6736 ( .A(\ImageBuffer[60][5] ), .B(\ImageBuffer[61][5] ), .C(
        \ImageBuffer[62][5] ), .D(\ImageBuffer[63][5] ), .S0(n3518), .S1(n3472), .Y(n4419) );
  MX4X1 U6737 ( .A(\ImageBuffer[44][5] ), .B(\ImageBuffer[45][5] ), .C(
        \ImageBuffer[46][5] ), .D(\ImageBuffer[47][5] ), .S0(n3522), .S1(n3474), .Y(n4424) );
  MX4X1 U6738 ( .A(\ImageBuffer[12][5] ), .B(\ImageBuffer[13][5] ), .C(
        \ImageBuffer[14][5] ), .D(\ImageBuffer[15][5] ), .S0(n3517), .S1(n3474), .Y(n4434) );
  MX4X1 U6739 ( .A(\ImageBuffer[60][6] ), .B(\ImageBuffer[61][6] ), .C(
        \ImageBuffer[62][6] ), .D(\ImageBuffer[63][6] ), .S0(n3518), .S1(n3474), .Y(n4439) );
  MX4X1 U6740 ( .A(\ImageBuffer[44][6] ), .B(\ImageBuffer[45][6] ), .C(
        \ImageBuffer[46][6] ), .D(\ImageBuffer[47][6] ), .S0(n3515), .S1(n3471), .Y(n4444) );
  MX4X1 U6741 ( .A(\ImageBuffer[12][6] ), .B(\ImageBuffer[13][6] ), .C(
        \ImageBuffer[14][6] ), .D(\ImageBuffer[15][6] ), .S0(n3512), .S1(n3472), .Y(n4454) );
  MX4X1 U6742 ( .A(\ImageBuffer[60][6] ), .B(\ImageBuffer[61][6] ), .C(
        \ImageBuffer[62][6] ), .D(\ImageBuffer[63][6] ), .S0(n3343), .S1(n3482), .Y(n4599) );
  MX4X1 U6743 ( .A(\ImageBuffer[44][6] ), .B(\ImageBuffer[45][6] ), .C(
        \ImageBuffer[46][6] ), .D(\ImageBuffer[47][6] ), .S0(n3506), .S1(n3484), .Y(n4604) );
  MX4X1 U6744 ( .A(\ImageBuffer[12][6] ), .B(\ImageBuffer[13][6] ), .C(
        \ImageBuffer[14][6] ), .D(\ImageBuffer[15][6] ), .S0(n3347), .S1(n3484), .Y(n4614) );
  MX4X1 U6745 ( .A(\ImageBuffer[60][7] ), .B(\ImageBuffer[61][7] ), .C(
        \ImageBuffer[62][7] ), .D(\ImageBuffer[63][7] ), .S0(n3515), .S1(n3473), .Y(n4459) );
  MX4X1 U6746 ( .A(\ImageBuffer[44][7] ), .B(\ImageBuffer[45][7] ), .C(
        \ImageBuffer[46][7] ), .D(\ImageBuffer[47][7] ), .S0(n3518), .S1(n3472), .Y(n4464) );
  MX4X1 U6747 ( .A(\ImageBuffer[12][7] ), .B(\ImageBuffer[13][7] ), .C(
        \ImageBuffer[14][7] ), .D(\ImageBuffer[15][7] ), .S0(n3521), .S1(n3471), .Y(n4474) );
  MX4X1 U6748 ( .A(\ImageBuffer[60][7] ), .B(\ImageBuffer[61][7] ), .C(
        \ImageBuffer[62][7] ), .D(\ImageBuffer[63][7] ), .S0(n3342), .S1(n3485), .Y(n4619) );
  MX4X1 U6749 ( .A(\ImageBuffer[44][7] ), .B(\ImageBuffer[45][7] ), .C(
        \ImageBuffer[46][7] ), .D(\ImageBuffer[47][7] ), .S0(n3506), .S1(n3482), .Y(n4624) );
  MX4X1 U6750 ( .A(\ImageBuffer[12][7] ), .B(\ImageBuffer[13][7] ), .C(
        \ImageBuffer[14][7] ), .D(\ImageBuffer[15][7] ), .S0(n3342), .S1(n3483), .Y(n4634) );
  MX4X1 U6751 ( .A(\ImageBuffer[44][4] ), .B(\ImageBuffer[45][4] ), .C(
        \ImageBuffer[46][4] ), .D(\ImageBuffer[47][4] ), .S0(n4119), .S1(n3749), .Y(n4033) );
  MX4X1 U6752 ( .A(\ImageBuffer[12][4] ), .B(\ImageBuffer[13][4] ), .C(
        \ImageBuffer[14][4] ), .D(\ImageBuffer[15][4] ), .S0(n3737), .S1(n3756), .Y(n4043) );
  MX4X1 U6753 ( .A(n4577), .B(n4575), .C(n4576), .D(n4574), .S0(n3496), .S1(
        n4640), .Y(n4578) );
  MX4X1 U6754 ( .A(\ImageBuffer[0][4] ), .B(\ImageBuffer[1][4] ), .C(
        \ImageBuffer[2][4] ), .D(\ImageBuffer[3][4] ), .S0(n3506), .S1(n3485), 
        .Y(n4577) );
  MX4X1 U6755 ( .A(\ImageBuffer[8][4] ), .B(\ImageBuffer[9][4] ), .C(
        \ImageBuffer[10][4] ), .D(\ImageBuffer[11][4] ), .S0(n3347), .S1(n3483), .Y(n4575) );
  MX4X1 U6756 ( .A(\ImageBuffer[12][4] ), .B(\ImageBuffer[13][4] ), .C(
        \ImageBuffer[14][4] ), .D(\ImageBuffer[15][4] ), .S0(n3343), .S1(n3483), .Y(n4574) );
  MX4X1 U6757 ( .A(n4597), .B(n4595), .C(n4596), .D(n4594), .S0(n3496), .S1(
        n4640), .Y(n4598) );
  MX4X1 U6758 ( .A(\ImageBuffer[0][5] ), .B(\ImageBuffer[1][5] ), .C(
        \ImageBuffer[2][5] ), .D(\ImageBuffer[3][5] ), .S0(n3343), .S1(n3482), 
        .Y(n4597) );
  MX4X1 U6759 ( .A(\ImageBuffer[8][5] ), .B(\ImageBuffer[9][5] ), .C(
        \ImageBuffer[10][5] ), .D(\ImageBuffer[11][5] ), .S0(n3506), .S1(n3485), .Y(n4595) );
  MX4X1 U6760 ( .A(\ImageBuffer[12][5] ), .B(\ImageBuffer[13][5] ), .C(
        \ImageBuffer[14][5] ), .D(\ImageBuffer[15][5] ), .S0(n3506), .S1(n3485), .Y(n4594) );
  MX4X1 U6761 ( .A(n3971), .B(n3969), .C(n3970), .D(n3968), .S0(n4109), .S1(
        n3758), .Y(n3972) );
  MX4X1 U6762 ( .A(\ImageBuffer[48][1] ), .B(\ImageBuffer[49][1] ), .C(
        \ImageBuffer[50][1] ), .D(\ImageBuffer[51][1] ), .S0(n3740), .S1(n3751), .Y(n3971) );
  MX4X1 U6763 ( .A(\ImageBuffer[56][1] ), .B(\ImageBuffer[57][1] ), .C(
        \ImageBuffer[58][1] ), .D(\ImageBuffer[59][1] ), .S0(n3735), .S1(n4125), .Y(n3969) );
  MX4X1 U6764 ( .A(\ImageBuffer[60][1] ), .B(\ImageBuffer[61][1] ), .C(
        \ImageBuffer[62][1] ), .D(\ImageBuffer[63][1] ), .S0(n4119), .S1(n4127), .Y(n3968) );
  MX4X1 U6765 ( .A(n4482), .B(n4480), .C(n4481), .D(n4479), .S0(n3496), .S1(
        n4641), .Y(n4483) );
  MX4X1 U6766 ( .A(\ImageBuffer[48][0] ), .B(\ImageBuffer[49][0] ), .C(
        \ImageBuffer[50][0] ), .D(\ImageBuffer[51][0] ), .S0(n3343), .S1(n3485), .Y(n4482) );
  MX4X1 U6767 ( .A(\ImageBuffer[56][0] ), .B(\ImageBuffer[57][0] ), .C(
        \ImageBuffer[58][0] ), .D(\ImageBuffer[59][0] ), .S0(n3347), .S1(n3484), .Y(n4480) );
  MX4X1 U6768 ( .A(\ImageBuffer[60][0] ), .B(\ImageBuffer[61][0] ), .C(
        \ImageBuffer[62][0] ), .D(\ImageBuffer[63][0] ), .S0(n3506), .S1(n3482), .Y(n4479) );
  MX4X1 U6769 ( .A(\ImageBuffer[48][1] ), .B(\ImageBuffer[49][1] ), .C(
        \ImageBuffer[50][1] ), .D(\ImageBuffer[51][1] ), .S0(n3516), .S1(n3474), .Y(n4342) );
  MX4X1 U6770 ( .A(\ImageBuffer[56][1] ), .B(\ImageBuffer[57][1] ), .C(
        \ImageBuffer[58][1] ), .D(\ImageBuffer[59][1] ), .S0(n3517), .S1(n3474), .Y(n4340) );
  MX4X1 U6771 ( .A(\ImageBuffer[48][2] ), .B(\ImageBuffer[49][2] ), .C(
        \ImageBuffer[50][2] ), .D(\ImageBuffer[51][2] ), .S0(n4115), .S1(n3753), .Y(n3991) );
  MX4X1 U6772 ( .A(\ImageBuffer[56][2] ), .B(\ImageBuffer[57][2] ), .C(
        \ImageBuffer[58][2] ), .D(\ImageBuffer[59][2] ), .S0(n4115), .S1(n4133), .Y(n3989) );
  MX4X1 U6773 ( .A(\ImageBuffer[60][2] ), .B(\ImageBuffer[61][2] ), .C(
        \ImageBuffer[62][2] ), .D(\ImageBuffer[63][2] ), .S0(n4115), .S1(n4132), .Y(n3988) );
  MX4X1 U6774 ( .A(\ImageBuffer[48][4] ), .B(\ImageBuffer[49][4] ), .C(
        \ImageBuffer[50][4] ), .D(\ImageBuffer[51][4] ), .S0(n3347), .S1(n3485), .Y(n4562) );
  MX4X1 U6775 ( .A(\ImageBuffer[56][4] ), .B(\ImageBuffer[57][4] ), .C(
        \ImageBuffer[58][4] ), .D(\ImageBuffer[59][4] ), .S0(n3347), .S1(n3483), .Y(n4560) );
  MX4X1 U6776 ( .A(\ImageBuffer[60][4] ), .B(\ImageBuffer[61][4] ), .C(
        \ImageBuffer[62][4] ), .D(\ImageBuffer[63][4] ), .S0(n3506), .S1(n3483), .Y(n4559) );
  MX4X1 U6777 ( .A(n4582), .B(n4580), .C(n4581), .D(n4579), .S0(n3496), .S1(
        n4640), .Y(n4583) );
  MX4X1 U6778 ( .A(\ImageBuffer[48][5] ), .B(\ImageBuffer[49][5] ), .C(
        \ImageBuffer[50][5] ), .D(\ImageBuffer[51][5] ), .S0(n3343), .S1(n3482), .Y(n4582) );
  MX4X1 U6779 ( .A(\ImageBuffer[56][5] ), .B(\ImageBuffer[57][5] ), .C(
        \ImageBuffer[58][5] ), .D(\ImageBuffer[59][5] ), .S0(n3506), .S1(n3482), .Y(n4580) );
  MX4X1 U6780 ( .A(\ImageBuffer[60][5] ), .B(\ImageBuffer[61][5] ), .C(
        \ImageBuffer[62][5] ), .D(\ImageBuffer[63][5] ), .S0(n3506), .S1(n3483), .Y(n4579) );
  MX4X1 U6781 ( .A(\ImageBuffer[48][2] ), .B(\ImageBuffer[49][2] ), .C(
        \ImageBuffer[50][2] ), .D(\ImageBuffer[51][2] ), .S0(n3486), .S1(n3924), .Y(n3803) );
  MX4X1 U6782 ( .A(\ImageBuffer[56][2] ), .B(\ImageBuffer[57][2] ), .C(
        \ImageBuffer[58][2] ), .D(\ImageBuffer[59][2] ), .S0(n5120), .S1(n3925), .Y(n3801) );
  MX4X1 U6783 ( .A(\ImageBuffer[60][2] ), .B(\ImageBuffer[61][2] ), .C(
        \ImageBuffer[62][2] ), .D(\ImageBuffer[63][2] ), .S0(n5120), .S1(n3921), .Y(n3800) );
  MX4X1 U6784 ( .A(n3616), .B(n3614), .C(n3615), .D(n3613), .S0(n3734), .S1(
        n3758), .Y(n3617) );
  MX4X1 U6785 ( .A(\ImageBuffer[48][2] ), .B(\ImageBuffer[49][2] ), .C(
        \ImageBuffer[50][2] ), .D(\ImageBuffer[51][2] ), .S0(n3745), .S1(n4126), .Y(n3616) );
  MX4X1 U6786 ( .A(\ImageBuffer[56][2] ), .B(\ImageBuffer[57][2] ), .C(
        \ImageBuffer[58][2] ), .D(\ImageBuffer[59][2] ), .S0(n3742), .S1(n3756), .Y(n3614) );
  MX4X1 U6787 ( .A(\ImageBuffer[60][2] ), .B(\ImageBuffer[61][2] ), .C(
        \ImageBuffer[62][2] ), .D(\ImageBuffer[63][2] ), .S0(n3743), .S1(n4125), .Y(n3613) );
  MX4X1 U6788 ( .A(\ImageBuffer[48][3] ), .B(\ImageBuffer[49][3] ), .C(
        \ImageBuffer[50][3] ), .D(\ImageBuffer[51][3] ), .S0(n3498), .S1(n4124), .Y(n3636) );
  MX4X1 U6789 ( .A(n4071), .B(n4069), .C(n4070), .D(n4068), .S0(n4109), .S1(
        n4136), .Y(n4072) );
  MX4X1 U6790 ( .A(\ImageBuffer[48][6] ), .B(\ImageBuffer[49][6] ), .C(
        \ImageBuffer[50][6] ), .D(\ImageBuffer[51][6] ), .S0(n4117), .S1(n3753), .Y(n4071) );
  MX4X1 U6791 ( .A(\ImageBuffer[56][6] ), .B(\ImageBuffer[57][6] ), .C(
        \ImageBuffer[58][6] ), .D(\ImageBuffer[59][6] ), .S0(n4117), .S1(n3753), .Y(n4069) );
  MX4X1 U6792 ( .A(\ImageBuffer[60][6] ), .B(\ImageBuffer[61][6] ), .C(
        \ImageBuffer[62][6] ), .D(\ImageBuffer[63][6] ), .S0(n4117), .S1(n4122), .Y(n4068) );
  MX4X1 U6793 ( .A(\ImageBuffer[48][3] ), .B(\ImageBuffer[49][3] ), .C(
        \ImageBuffer[50][3] ), .D(\ImageBuffer[51][3] ), .S0(n4116), .S1(n4126), .Y(n4011) );
  MX4X1 U6794 ( .A(\ImageBuffer[48][4] ), .B(\ImageBuffer[49][4] ), .C(
        \ImageBuffer[50][4] ), .D(\ImageBuffer[51][4] ), .S0(n3742), .S1(n4130), .Y(n3656) );
  MX4X1 U6795 ( .A(\ImageBuffer[56][4] ), .B(\ImageBuffer[57][4] ), .C(
        \ImageBuffer[58][4] ), .D(\ImageBuffer[59][4] ), .S0(n3742), .S1(n3755), .Y(n3654) );
  MX4X1 U6796 ( .A(\ImageBuffer[60][4] ), .B(\ImageBuffer[61][4] ), .C(
        \ImageBuffer[62][4] ), .D(\ImageBuffer[63][4] ), .S0(n3742), .S1(n4134), .Y(n3653) );
  MX4X1 U6797 ( .A(n4542), .B(n4540), .C(n4541), .D(n4539), .S0(n3496), .S1(
        n4639), .Y(n4543) );
  MX4X1 U6798 ( .A(\ImageBuffer[48][3] ), .B(\ImageBuffer[49][3] ), .C(
        \ImageBuffer[50][3] ), .D(\ImageBuffer[51][3] ), .S0(n3343), .S1(n3484), .Y(n4542) );
  MX4X1 U6799 ( .A(\ImageBuffer[52][3] ), .B(\ImageBuffer[53][3] ), .C(
        \ImageBuffer[54][3] ), .D(\ImageBuffer[55][3] ), .S0(n3343), .S1(n3485), .Y(n4541) );
  MX4X1 U6800 ( .A(n4031), .B(n4029), .C(n4030), .D(n4028), .S0(n4108), .S1(
        n4135), .Y(n4032) );
  MX4X1 U6801 ( .A(\ImageBuffer[48][4] ), .B(\ImageBuffer[49][4] ), .C(
        \ImageBuffer[50][4] ), .D(\ImageBuffer[51][4] ), .S0(n4119), .S1(n3753), .Y(n4031) );
  MX4X1 U6802 ( .A(\ImageBuffer[56][4] ), .B(\ImageBuffer[57][4] ), .C(
        \ImageBuffer[58][4] ), .D(\ImageBuffer[59][4] ), .S0(n4119), .S1(n3748), .Y(n4029) );
  MX4X1 U6803 ( .A(\ImageBuffer[60][4] ), .B(\ImageBuffer[61][4] ), .C(
        \ImageBuffer[62][4] ), .D(\ImageBuffer[63][4] ), .S0(n4119), .S1(n3756), .Y(n4028) );
  MX4X1 U6804 ( .A(\ImageBuffer[40][2] ), .B(\ImageBuffer[41][2] ), .C(
        \ImageBuffer[42][2] ), .D(\ImageBuffer[43][2] ), .S0(n3740), .S1(n3754), .Y(n3994) );
  MX4X1 U6805 ( .A(\ImageBuffer[8][2] ), .B(\ImageBuffer[9][2] ), .C(
        \ImageBuffer[10][2] ), .D(\ImageBuffer[11][2] ), .S0(n3735), .S1(n3754), .Y(n4004) );
  MX4X1 U6806 ( .A(\ImageBuffer[56][0] ), .B(\ImageBuffer[57][0] ), .C(
        \ImageBuffer[58][0] ), .D(\ImageBuffer[59][0] ), .S0(n4114), .S1(n3757), .Y(n3951) );
  MX4X1 U6807 ( .A(\ImageBuffer[40][2] ), .B(\ImageBuffer[41][2] ), .C(
        \ImageBuffer[42][2] ), .D(\ImageBuffer[43][2] ), .S0(n3939), .S1(n3923), .Y(n3806) );
  MX4X1 U6808 ( .A(\ImageBuffer[8][2] ), .B(\ImageBuffer[9][2] ), .C(
        \ImageBuffer[10][2] ), .D(\ImageBuffer[11][2] ), .S0(n3939), .S1(n3925), .Y(n3816) );
  MX4X1 U6809 ( .A(\ImageBuffer[56][0] ), .B(\ImageBuffer[57][0] ), .C(
        \ImageBuffer[58][0] ), .D(\ImageBuffer[59][0] ), .S0(n4117), .S1(n3750), .Y(n3574) );
  MX4X1 U6810 ( .A(\ImageBuffer[40][0] ), .B(\ImageBuffer[41][0] ), .C(
        \ImageBuffer[42][0] ), .D(\ImageBuffer[43][0] ), .S0(n4119), .S1(n3756), .Y(n3579) );
  MX4X1 U6811 ( .A(\ImageBuffer[56][0] ), .B(\ImageBuffer[57][0] ), .C(
        \ImageBuffer[58][0] ), .D(\ImageBuffer[59][0] ), .S0(n3938), .S1(n3929), .Y(n3761) );
  MX4X1 U6812 ( .A(\ImageBuffer[40][0] ), .B(\ImageBuffer[41][0] ), .C(
        \ImageBuffer[42][0] ), .D(\ImageBuffer[43][0] ), .S0(n3938), .S1(n5123), .Y(n3766) );
  MX4X1 U6813 ( .A(\ImageBuffer[56][2] ), .B(\ImageBuffer[57][2] ), .C(
        \ImageBuffer[58][2] ), .D(\ImageBuffer[59][2] ), .S0(n3506), .S1(n3483), .Y(n4520) );
  MX4X1 U6814 ( .A(\ImageBuffer[8][2] ), .B(\ImageBuffer[9][2] ), .C(
        \ImageBuffer[10][2] ), .D(\ImageBuffer[11][2] ), .S0(n3506), .S1(n3483), .Y(n4535) );
  MX4X1 U6815 ( .A(\ImageBuffer[40][2] ), .B(\ImageBuffer[41][2] ), .C(
        \ImageBuffer[42][2] ), .D(\ImageBuffer[43][2] ), .S0(n3741), .S1(n4125), .Y(n3619) );
  MX4X1 U6816 ( .A(\ImageBuffer[8][2] ), .B(\ImageBuffer[9][2] ), .C(
        \ImageBuffer[10][2] ), .D(\ImageBuffer[11][2] ), .S0(n3741), .S1(n3748), .Y(n3629) );
  MX4X1 U6817 ( .A(\ImageBuffer[40][3] ), .B(\ImageBuffer[41][3] ), .C(
        \ImageBuffer[42][3] ), .D(\ImageBuffer[43][3] ), .S0(n3498), .S1(n4126), .Y(n3639) );
  MX4X1 U6818 ( .A(\ImageBuffer[8][3] ), .B(\ImageBuffer[9][3] ), .C(
        \ImageBuffer[10][3] ), .D(\ImageBuffer[11][3] ), .S0(n3498), .S1(n4130), .Y(n3649) );
  MX4X1 U6819 ( .A(\ImageBuffer[24][6] ), .B(\ImageBuffer[25][6] ), .C(
        \ImageBuffer[26][6] ), .D(\ImageBuffer[27][6] ), .S0(n3488), .S1(n3750), .Y(n3704) );
  MX4X1 U6820 ( .A(\ImageBuffer[56][6] ), .B(\ImageBuffer[57][6] ), .C(
        \ImageBuffer[58][6] ), .D(\ImageBuffer[59][6] ), .S0(n3743), .S1(n3748), .Y(n3694) );
  MX4X1 U6821 ( .A(\ImageBuffer[8][5] ), .B(\ImageBuffer[9][5] ), .C(
        \ImageBuffer[10][5] ), .D(\ImageBuffer[11][5] ), .S0(n4117), .S1(n4134), .Y(n4064) );
  MX4X1 U6822 ( .A(\ImageBuffer[8][6] ), .B(\ImageBuffer[9][6] ), .C(
        \ImageBuffer[10][6] ), .D(\ImageBuffer[11][6] ), .S0(n4118), .S1(n3756), .Y(n4084) );
  MX4X1 U6823 ( .A(\ImageBuffer[8][3] ), .B(\ImageBuffer[9][3] ), .C(
        \ImageBuffer[10][3] ), .D(\ImageBuffer[11][3] ), .S0(n4116), .S1(n3752), .Y(n4024) );
  MX4X1 U6824 ( .A(\ImageBuffer[40][3] ), .B(\ImageBuffer[41][3] ), .C(
        \ImageBuffer[42][3] ), .D(\ImageBuffer[43][3] ), .S0(n3489), .S1(n3924), .Y(n3826) );
  MX4X1 U6825 ( .A(\ImageBuffer[40][4] ), .B(\ImageBuffer[41][4] ), .C(
        \ImageBuffer[42][4] ), .D(\ImageBuffer[43][4] ), .S0(n3742), .S1(n4125), .Y(n3659) );
  MX4X1 U6826 ( .A(\ImageBuffer[8][4] ), .B(\ImageBuffer[9][4] ), .C(
        \ImageBuffer[10][4] ), .D(\ImageBuffer[11][4] ), .S0(n3498), .S1(n4126), .Y(n3669) );
  MX4X1 U6827 ( .A(\ImageBuffer[40][4] ), .B(\ImageBuffer[41][4] ), .C(
        \ImageBuffer[42][4] ), .D(\ImageBuffer[43][4] ), .S0(n3486), .S1(n3922), .Y(n3846) );
  MX4X1 U6828 ( .A(\ImageBuffer[8][4] ), .B(\ImageBuffer[9][4] ), .C(
        \ImageBuffer[10][4] ), .D(\ImageBuffer[11][4] ), .S0(n3939), .S1(n3931), .Y(n3856) );
  MX4X1 U6829 ( .A(\ImageBuffer[56][2] ), .B(\ImageBuffer[57][2] ), .C(
        \ImageBuffer[58][2] ), .D(\ImageBuffer[59][2] ), .S0(n4300), .S1(n5113), .Y(n4178) );
  MX4X1 U6830 ( .A(\ImageBuffer[8][2] ), .B(\ImageBuffer[9][2] ), .C(
        \ImageBuffer[10][2] ), .D(\ImageBuffer[11][2] ), .S0(n3938), .S1(n4314), .Y(n4193) );
  MX4X1 U6831 ( .A(\ImageBuffer[40][2] ), .B(\ImageBuffer[41][2] ), .C(
        \ImageBuffer[42][2] ), .D(\ImageBuffer[43][2] ), .S0(n3938), .S1(n4304), .Y(n4183) );
  MX4X1 U6832 ( .A(\ImageBuffer[40][6] ), .B(\ImageBuffer[41][6] ), .C(
        \ImageBuffer[42][6] ), .D(\ImageBuffer[43][6] ), .S0(n4300), .S1(n3341), .Y(n3886) );
  MX4X1 U6833 ( .A(\ImageBuffer[8][6] ), .B(\ImageBuffer[9][6] ), .C(
        \ImageBuffer[10][6] ), .D(\ImageBuffer[11][6] ), .S0(n3935), .S1(n3920), .Y(n3896) );
  MX4X1 U6834 ( .A(\ImageBuffer[40][4] ), .B(\ImageBuffer[41][4] ), .C(
        \ImageBuffer[42][4] ), .D(\ImageBuffer[43][4] ), .S0(n3940), .S1(n4306), .Y(n4223) );
  MX4X1 U6835 ( .A(\ImageBuffer[24][4] ), .B(\ImageBuffer[25][4] ), .C(
        \ImageBuffer[26][4] ), .D(\ImageBuffer[27][4] ), .S0(n3935), .S1(n4312), .Y(n4228) );
  MX4X1 U6836 ( .A(\ImageBuffer[56][4] ), .B(\ImageBuffer[57][4] ), .C(
        \ImageBuffer[58][4] ), .D(\ImageBuffer[59][4] ), .S0(n3941), .S1(n4317), .Y(n4218) );
  MX4X1 U6837 ( .A(\ImageBuffer[8][6] ), .B(\ImageBuffer[9][6] ), .C(
        \ImageBuffer[10][6] ), .D(\ImageBuffer[11][6] ), .S0(n4297), .S1(n4313), .Y(n4273) );
  MX4X1 U6838 ( .A(\ImageBuffer[56][0] ), .B(\ImageBuffer[57][0] ), .C(
        \ImageBuffer[58][0] ), .D(\ImageBuffer[59][0] ), .S0(n3939), .S1(n4316), .Y(n4138) );
  MX4X1 U6839 ( .A(\ImageBuffer[8][0] ), .B(\ImageBuffer[9][0] ), .C(
        \ImageBuffer[10][0] ), .D(\ImageBuffer[11][0] ), .S0(n3939), .S1(n4317), .Y(n4153) );
  MX4X1 U6840 ( .A(\ImageBuffer[40][0] ), .B(\ImageBuffer[41][0] ), .C(
        \ImageBuffer[42][0] ), .D(\ImageBuffer[43][0] ), .S0(n3938), .S1(n4311), .Y(n4143) );
  MX4X1 U6841 ( .A(\ImageBuffer[24][0] ), .B(\ImageBuffer[25][0] ), .C(
        \ImageBuffer[26][0] ), .D(\ImageBuffer[27][0] ), .S0(n3511), .S1(n3471), .Y(n4330) );
  MX4X1 U6842 ( .A(\ImageBuffer[8][0] ), .B(\ImageBuffer[9][0] ), .C(
        \ImageBuffer[10][0] ), .D(\ImageBuffer[11][0] ), .S0(n3513), .S1(n3471), .Y(n4335) );
  MX4X1 U6843 ( .A(\ImageBuffer[40][0] ), .B(\ImageBuffer[41][0] ), .C(
        \ImageBuffer[42][0] ), .D(\ImageBuffer[43][0] ), .S0(n3513), .S1(n3471), .Y(n4325) );
  MX4X1 U6844 ( .A(\ImageBuffer[24][1] ), .B(\ImageBuffer[25][1] ), .C(
        \ImageBuffer[26][1] ), .D(\ImageBuffer[27][1] ), .S0(n3506), .S1(n3483), .Y(n4510) );
  MX4X1 U6845 ( .A(\ImageBuffer[40][1] ), .B(\ImageBuffer[41][1] ), .C(
        \ImageBuffer[42][1] ), .D(\ImageBuffer[43][1] ), .S0(n3343), .S1(n3483), .Y(n4505) );
  MX4X1 U6846 ( .A(\ImageBuffer[8][1] ), .B(\ImageBuffer[9][1] ), .C(
        \ImageBuffer[10][1] ), .D(\ImageBuffer[11][1] ), .S0(n3347), .S1(n3484), .Y(n4515) );
  MX4X1 U6847 ( .A(\ImageBuffer[24][3] ), .B(\ImageBuffer[25][3] ), .C(
        \ImageBuffer[26][3] ), .D(\ImageBuffer[27][3] ), .S0(n3511), .S1(n3474), .Y(n4390) );
  MX4X1 U6848 ( .A(\ImageBuffer[40][3] ), .B(\ImageBuffer[41][3] ), .C(
        \ImageBuffer[42][3] ), .D(\ImageBuffer[43][3] ), .S0(n3514), .S1(n3473), .Y(n4385) );
  MX4X1 U6849 ( .A(\ImageBuffer[8][3] ), .B(\ImageBuffer[9][3] ), .C(
        \ImageBuffer[10][3] ), .D(\ImageBuffer[11][3] ), .S0(n3512), .S1(n3471), .Y(n4395) );
  MX4X1 U6850 ( .A(\ImageBuffer[56][4] ), .B(\ImageBuffer[57][4] ), .C(
        \ImageBuffer[58][4] ), .D(\ImageBuffer[59][4] ), .S0(n3519), .S1(n3472), .Y(n4400) );
  MX4X1 U6851 ( .A(\ImageBuffer[40][4] ), .B(\ImageBuffer[41][4] ), .C(
        \ImageBuffer[42][4] ), .D(\ImageBuffer[43][4] ), .S0(n3514), .S1(n3473), .Y(n4405) );
  MX4X1 U6852 ( .A(\ImageBuffer[8][4] ), .B(\ImageBuffer[9][4] ), .C(
        \ImageBuffer[10][4] ), .D(\ImageBuffer[11][4] ), .S0(n3515), .S1(n3473), .Y(n4415) );
  MX4X1 U6853 ( .A(\ImageBuffer[56][5] ), .B(\ImageBuffer[57][5] ), .C(
        \ImageBuffer[58][5] ), .D(\ImageBuffer[59][5] ), .S0(n3514), .S1(n3474), .Y(n4420) );
  MX4X1 U6854 ( .A(\ImageBuffer[40][5] ), .B(\ImageBuffer[41][5] ), .C(
        \ImageBuffer[42][5] ), .D(\ImageBuffer[43][5] ), .S0(n3516), .S1(n3471), .Y(n4425) );
  MX4X1 U6855 ( .A(\ImageBuffer[8][5] ), .B(\ImageBuffer[9][5] ), .C(
        \ImageBuffer[10][5] ), .D(\ImageBuffer[11][5] ), .S0(n3518), .S1(n3472), .Y(n4435) );
  MX4X1 U6856 ( .A(\ImageBuffer[56][6] ), .B(\ImageBuffer[57][6] ), .C(
        \ImageBuffer[58][6] ), .D(\ImageBuffer[59][6] ), .S0(n3514), .S1(n3474), .Y(n4440) );
  MX4X1 U6857 ( .A(\ImageBuffer[40][6] ), .B(\ImageBuffer[41][6] ), .C(
        \ImageBuffer[42][6] ), .D(\ImageBuffer[43][6] ), .S0(n3515), .S1(n3472), .Y(n4445) );
  MX4X1 U6858 ( .A(\ImageBuffer[8][6] ), .B(\ImageBuffer[9][6] ), .C(
        \ImageBuffer[10][6] ), .D(\ImageBuffer[11][6] ), .S0(n3511), .S1(n3474), .Y(n4455) );
  MX4X1 U6859 ( .A(\ImageBuffer[56][6] ), .B(\ImageBuffer[57][6] ), .C(
        \ImageBuffer[58][6] ), .D(\ImageBuffer[59][6] ), .S0(n3343), .S1(n3483), .Y(n4600) );
  MX4X1 U6860 ( .A(\ImageBuffer[40][6] ), .B(\ImageBuffer[41][6] ), .C(
        \ImageBuffer[42][6] ), .D(\ImageBuffer[43][6] ), .S0(n3347), .S1(n3482), .Y(n4605) );
  MX4X1 U6861 ( .A(\ImageBuffer[8][6] ), .B(\ImageBuffer[9][6] ), .C(
        \ImageBuffer[10][6] ), .D(\ImageBuffer[11][6] ), .S0(n3343), .S1(n3485), .Y(n4615) );
  MX4X1 U6862 ( .A(\ImageBuffer[56][7] ), .B(\ImageBuffer[57][7] ), .C(
        \ImageBuffer[58][7] ), .D(\ImageBuffer[59][7] ), .S0(n3517), .S1(n3474), .Y(n4460) );
  MX4X1 U6863 ( .A(\ImageBuffer[40][7] ), .B(\ImageBuffer[41][7] ), .C(
        \ImageBuffer[42][7] ), .D(\ImageBuffer[43][7] ), .S0(n3514), .S1(n3471), .Y(n4465) );
  MX4X1 U6864 ( .A(\ImageBuffer[8][7] ), .B(\ImageBuffer[9][7] ), .C(
        \ImageBuffer[10][7] ), .D(\ImageBuffer[11][7] ), .S0(n3511), .S1(n3471), .Y(n4475) );
  MX4X1 U6865 ( .A(\ImageBuffer[56][7] ), .B(\ImageBuffer[57][7] ), .C(
        \ImageBuffer[58][7] ), .D(\ImageBuffer[59][7] ), .S0(n3342), .S1(n3485), .Y(n4620) );
  MX4X1 U6866 ( .A(\ImageBuffer[40][7] ), .B(\ImageBuffer[41][7] ), .C(
        \ImageBuffer[42][7] ), .D(\ImageBuffer[43][7] ), .S0(n3506), .S1(n3485), .Y(n4625) );
  MX4X1 U6867 ( .A(\ImageBuffer[8][7] ), .B(\ImageBuffer[9][7] ), .C(
        \ImageBuffer[10][7] ), .D(\ImageBuffer[11][7] ), .S0(n3346), .S1(n3483), .Y(n4635) );
  MX4X1 U6868 ( .A(\ImageBuffer[40][4] ), .B(\ImageBuffer[41][4] ), .C(
        \ImageBuffer[42][4] ), .D(\ImageBuffer[43][4] ), .S0(n4119), .S1(N2494), .Y(n4034) );
  MX4X1 U6869 ( .A(\ImageBuffer[8][4] ), .B(\ImageBuffer[9][4] ), .C(
        \ImageBuffer[10][4] ), .D(\ImageBuffer[11][4] ), .S0(n4116), .S1(n3756), .Y(n4044) );
  MX4X1 U6870 ( .A(n4567), .B(n4565), .C(n4566), .D(n4564), .S0(n3496), .S1(
        n4639), .Y(n4568) );
  MX4X1 U6871 ( .A(\ImageBuffer[32][4] ), .B(\ImageBuffer[33][4] ), .C(
        \ImageBuffer[34][4] ), .D(\ImageBuffer[35][4] ), .S0(n3506), .S1(n3482), .Y(n4567) );
  MX4X1 U6872 ( .A(\ImageBuffer[40][4] ), .B(\ImageBuffer[41][4] ), .C(
        \ImageBuffer[42][4] ), .D(\ImageBuffer[43][4] ), .S0(n3506), .S1(n3484), .Y(n4565) );
  MX4X1 U6873 ( .A(\ImageBuffer[44][4] ), .B(\ImageBuffer[45][4] ), .C(
        \ImageBuffer[46][4] ), .D(\ImageBuffer[47][4] ), .S0(n3347), .S1(n3482), .Y(n4564) );
  MX4X1 U6874 ( .A(n4587), .B(n4585), .C(n4586), .D(n4584), .S0(n3496), .S1(
        n4640), .Y(n4588) );
  MX4X1 U6875 ( .A(\ImageBuffer[32][5] ), .B(\ImageBuffer[33][5] ), .C(
        \ImageBuffer[34][5] ), .D(\ImageBuffer[35][5] ), .S0(n3506), .S1(n3483), .Y(n4587) );
  MX4X1 U6876 ( .A(\ImageBuffer[40][5] ), .B(\ImageBuffer[41][5] ), .C(
        \ImageBuffer[42][5] ), .D(\ImageBuffer[43][5] ), .S0(n3347), .S1(n3484), .Y(n4585) );
  MX4X1 U6877 ( .A(\ImageBuffer[44][5] ), .B(\ImageBuffer[45][5] ), .C(
        \ImageBuffer[46][5] ), .D(\ImageBuffer[47][5] ), .S0(n3343), .S1(n3482), .Y(n4584) );
  MX4X1 U6878 ( .A(n3976), .B(n3974), .C(n3975), .D(n3973), .S0(n4109), .S1(
        n3758), .Y(n3977) );
  MX4X1 U6879 ( .A(\ImageBuffer[32][1] ), .B(\ImageBuffer[33][1] ), .C(
        \ImageBuffer[34][1] ), .D(\ImageBuffer[35][1] ), .S0(n3735), .S1(n3755), .Y(n3976) );
  MX4X1 U6880 ( .A(\ImageBuffer[40][1] ), .B(\ImageBuffer[41][1] ), .C(
        \ImageBuffer[42][1] ), .D(\ImageBuffer[43][1] ), .S0(n3740), .S1(n4126), .Y(n3974) );
  MX4X1 U6881 ( .A(\ImageBuffer[44][1] ), .B(\ImageBuffer[45][1] ), .C(
        \ImageBuffer[46][1] ), .D(\ImageBuffer[47][1] ), .S0(n3735), .S1(N2494), .Y(n3973) );
  MX4X1 U6882 ( .A(n4487), .B(n4485), .C(n4486), .D(n4484), .S0(n3496), .S1(
        n4641), .Y(n4488) );
  MX4X1 U6883 ( .A(\ImageBuffer[32][0] ), .B(\ImageBuffer[33][0] ), .C(
        \ImageBuffer[34][0] ), .D(\ImageBuffer[35][0] ), .S0(n3347), .S1(n3484), .Y(n4487) );
  MX4X1 U6884 ( .A(\ImageBuffer[40][0] ), .B(\ImageBuffer[41][0] ), .C(
        \ImageBuffer[42][0] ), .D(\ImageBuffer[43][0] ), .S0(n3506), .S1(n3482), .Y(n4485) );
  MX4X1 U6885 ( .A(\ImageBuffer[44][0] ), .B(\ImageBuffer[45][0] ), .C(
        \ImageBuffer[46][0] ), .D(\ImageBuffer[47][0] ), .S0(n3506), .S1(n3484), .Y(n4484) );
  MX4X1 U6886 ( .A(n4347), .B(n4345), .C(n4346), .D(n4344), .S0(n3503), .S1(
        n3495), .Y(n4348) );
  MX4X1 U6887 ( .A(\ImageBuffer[32][1] ), .B(\ImageBuffer[33][1] ), .C(
        \ImageBuffer[34][1] ), .D(\ImageBuffer[35][1] ), .S0(n3511), .S1(n3471), .Y(n4347) );
  MX4X1 U6888 ( .A(\ImageBuffer[40][1] ), .B(\ImageBuffer[41][1] ), .C(
        \ImageBuffer[42][1] ), .D(\ImageBuffer[43][1] ), .S0(n3513), .S1(n3471), .Y(n4345) );
  MX4X1 U6889 ( .A(\ImageBuffer[44][1] ), .B(\ImageBuffer[45][1] ), .C(
        \ImageBuffer[46][1] ), .D(\ImageBuffer[47][1] ), .S0(n3512), .S1(n3472), .Y(n4344) );
  MX4X1 U6890 ( .A(n3701), .B(n3699), .C(n3700), .D(n3698), .S0(n3734), .S1(
        n3759), .Y(n3702) );
  MX4X1 U6891 ( .A(\ImageBuffer[44][6] ), .B(\ImageBuffer[45][6] ), .C(
        \ImageBuffer[46][6] ), .D(\ImageBuffer[47][6] ), .S0(n3743), .S1(n3754), .Y(n3698) );
  MX4X1 U6892 ( .A(\ImageBuffer[36][6] ), .B(\ImageBuffer[37][6] ), .C(
        \ImageBuffer[38][6] ), .D(\ImageBuffer[39][6] ), .S0(n4115), .S1(n4124), .Y(n3700) );
  MX4X1 U6893 ( .A(\ImageBuffer[40][6] ), .B(\ImageBuffer[41][6] ), .C(
        \ImageBuffer[42][6] ), .D(\ImageBuffer[43][6] ), .S0(n3743), .S1(n3750), .Y(n3699) );
  MX4X1 U6894 ( .A(n4076), .B(n4074), .C(n4075), .D(n4073), .S0(n4109), .S1(
        n4136), .Y(n4077) );
  MX4X1 U6895 ( .A(\ImageBuffer[32][6] ), .B(\ImageBuffer[33][6] ), .C(
        \ImageBuffer[34][6] ), .D(\ImageBuffer[35][6] ), .S0(n4118), .S1(n3752), .Y(n4076) );
  MX4X1 U6896 ( .A(\ImageBuffer[40][6] ), .B(\ImageBuffer[41][6] ), .C(
        \ImageBuffer[42][6] ), .D(\ImageBuffer[43][6] ), .S0(n4117), .S1(n4127), .Y(n4074) );
  MX4X1 U6897 ( .A(\ImageBuffer[44][6] ), .B(\ImageBuffer[45][6] ), .C(
        \ImageBuffer[46][6] ), .D(\ImageBuffer[47][6] ), .S0(n4117), .S1(n3755), .Y(n4073) );
  MX4X1 U6898 ( .A(\ImageBuffer[32][3] ), .B(\ImageBuffer[33][3] ), .C(
        \ImageBuffer[34][3] ), .D(\ImageBuffer[35][3] ), .S0(n4116), .S1(n3749), .Y(n4016) );
  MX4X1 U6899 ( .A(\ImageBuffer[40][3] ), .B(\ImageBuffer[41][3] ), .C(
        \ImageBuffer[42][3] ), .D(\ImageBuffer[43][3] ), .S0(n4116), .S1(n4122), .Y(n4014) );
  MX4X1 U6900 ( .A(\ImageBuffer[44][3] ), .B(\ImageBuffer[45][3] ), .C(
        \ImageBuffer[46][3] ), .D(\ImageBuffer[47][3] ), .S0(n4116), .S1(n4124), .Y(n4013) );
  MX4X1 U6901 ( .A(n4547), .B(n4545), .C(n4546), .D(n4544), .S0(n3496), .S1(
        n4639), .Y(n4548) );
  MX4X1 U6902 ( .A(\ImageBuffer[32][3] ), .B(\ImageBuffer[33][3] ), .C(
        \ImageBuffer[34][3] ), .D(\ImageBuffer[35][3] ), .S0(n3506), .S1(n3483), .Y(n4547) );
  MX4X1 U6903 ( .A(\ImageBuffer[40][3] ), .B(\ImageBuffer[41][3] ), .C(
        \ImageBuffer[42][3] ), .D(\ImageBuffer[43][3] ), .S0(n3347), .S1(n3484), .Y(n4545) );
  MX4X1 U6904 ( .A(\ImageBuffer[44][3] ), .B(\ImageBuffer[45][3] ), .C(
        \ImageBuffer[46][3] ), .D(\ImageBuffer[47][3] ), .S0(n3347), .S1(n3485), .Y(n4544) );
  MX4X1 U6905 ( .A(n4382), .B(n4380), .C(n4381), .D(n4379), .S0(n3503), .S1(
        n3495), .Y(n4383) );
  MX4X1 U6906 ( .A(\ImageBuffer[48][3] ), .B(\ImageBuffer[49][3] ), .C(
        \ImageBuffer[50][3] ), .D(\ImageBuffer[51][3] ), .S0(n3522), .S1(n3472), .Y(n4382) );
  MX4X1 U6907 ( .A(\ImageBuffer[56][3] ), .B(\ImageBuffer[57][3] ), .C(
        \ImageBuffer[58][3] ), .D(\ImageBuffer[59][3] ), .S0(n3513), .S1(n3472), .Y(n4380) );
  MX4X1 U6908 ( .A(\ImageBuffer[60][3] ), .B(\ImageBuffer[61][3] ), .C(
        \ImageBuffer[62][3] ), .D(\ImageBuffer[63][3] ), .S0(n3511), .S1(n3474), .Y(n4379) );
  MX4X1 U6909 ( .A(n4322), .B(n4320), .C(n4321), .D(n4319), .S0(n3503), .S1(
        n3495), .Y(n4323) );
  MX4X1 U6910 ( .A(\ImageBuffer[48][0] ), .B(\ImageBuffer[49][0] ), .C(
        \ImageBuffer[50][0] ), .D(\ImageBuffer[51][0] ), .S0(n3517), .S1(n3474), .Y(n4322) );
  MX4X1 U6911 ( .A(\ImageBuffer[56][0] ), .B(\ImageBuffer[57][0] ), .C(
        \ImageBuffer[58][0] ), .D(\ImageBuffer[59][0] ), .S0(n3516), .S1(n3473), .Y(n4320) );
  MX4X1 U6912 ( .A(\ImageBuffer[60][0] ), .B(\ImageBuffer[61][0] ), .C(
        \ImageBuffer[62][0] ), .D(\ImageBuffer[63][0] ), .S0(n3517), .S1(n3471), .Y(n4319) );
  MX4X1 U6913 ( .A(n3843), .B(n3841), .C(n3842), .D(n3840), .S0(n3933), .S1(
        n3409), .Y(n3844) );
  MX4X1 U6914 ( .A(\ImageBuffer[60][4] ), .B(\ImageBuffer[61][4] ), .C(
        \ImageBuffer[62][4] ), .D(\ImageBuffer[63][4] ), .S0(n3486), .S1(n3932), .Y(n3840) );
  MX4X1 U6915 ( .A(\ImageBuffer[52][4] ), .B(\ImageBuffer[53][4] ), .C(
        \ImageBuffer[54][4] ), .D(\ImageBuffer[55][4] ), .S0(n3486), .S1(n3340), .Y(n3842) );
  MX4X1 U6916 ( .A(\ImageBuffer[56][4] ), .B(\ImageBuffer[57][4] ), .C(
        \ImageBuffer[58][4] ), .D(\ImageBuffer[59][4] ), .S0(n3486), .S1(n3931), .Y(n3841) );
  MX4X1 U6917 ( .A(\ImageBuffer[48][1] ), .B(\ImageBuffer[49][1] ), .C(
        \ImageBuffer[50][1] ), .D(\ImageBuffer[51][1] ), .S0(n3939), .S1(n3926), .Y(n3783) );
  MX4X1 U6918 ( .A(\ImageBuffer[56][1] ), .B(\ImageBuffer[57][1] ), .C(
        \ImageBuffer[58][1] ), .D(\ImageBuffer[59][1] ), .S0(n3939), .S1(n3931), .Y(n3781) );
  MX4X1 U6919 ( .A(\ImageBuffer[60][1] ), .B(\ImageBuffer[61][1] ), .C(
        \ImageBuffer[62][1] ), .D(\ImageBuffer[63][1] ), .S0(n3939), .S1(n3930), .Y(n3780) );
  MX4X1 U6920 ( .A(n4502), .B(n4500), .C(n4501), .D(n4499), .S0(n3496), .S1(
        n4641), .Y(n4503) );
  MX4X1 U6921 ( .A(\ImageBuffer[48][1] ), .B(\ImageBuffer[49][1] ), .C(
        \ImageBuffer[50][1] ), .D(\ImageBuffer[51][1] ), .S0(n3506), .S1(n3485), .Y(n4502) );
  MX4X1 U6922 ( .A(\ImageBuffer[56][1] ), .B(\ImageBuffer[57][1] ), .C(
        \ImageBuffer[58][1] ), .D(\ImageBuffer[59][1] ), .S0(n3506), .S1(n3484), .Y(n4500) );
  MX4X1 U6923 ( .A(\ImageBuffer[60][1] ), .B(\ImageBuffer[61][1] ), .C(
        \ImageBuffer[62][1] ), .D(\ImageBuffer[63][1] ), .S0(n3347), .S1(n3485), .Y(n4499) );
  MX4X1 U6924 ( .A(n3838), .B(n3836), .C(n3837), .D(n3835), .S0(n3933), .S1(
        n3409), .Y(n3839) );
  MX4X1 U6925 ( .A(\ImageBuffer[12][3] ), .B(\ImageBuffer[13][3] ), .C(
        \ImageBuffer[14][3] ), .D(\ImageBuffer[15][3] ), .S0(n3489), .S1(n3480), .Y(n3835) );
  MX4X1 U6926 ( .A(\ImageBuffer[4][3] ), .B(\ImageBuffer[5][3] ), .C(
        \ImageBuffer[6][3] ), .D(\ImageBuffer[7][3] ), .S0(n3489), .S1(n3920), 
        .Y(n3837) );
  MX4X1 U6927 ( .A(\ImageBuffer[8][3] ), .B(\ImageBuffer[9][3] ), .C(
        \ImageBuffer[10][3] ), .D(\ImageBuffer[11][3] ), .S0(n3489), .S1(n3340), .Y(n3836) );
  MX4X1 U6928 ( .A(n3833), .B(n3831), .C(n3832), .D(n3830), .S0(n3933), .S1(
        n3409), .Y(n3834) );
  MX4X1 U6929 ( .A(\ImageBuffer[28][3] ), .B(\ImageBuffer[29][3] ), .C(
        \ImageBuffer[30][3] ), .D(\ImageBuffer[31][3] ), .S0(n3489), .S1(n3921), .Y(n3830) );
  MX4X1 U6930 ( .A(\ImageBuffer[20][3] ), .B(\ImageBuffer[21][3] ), .C(
        \ImageBuffer[22][3] ), .D(\ImageBuffer[23][3] ), .S0(n3489), .S1(n3932), .Y(n3832) );
  MX4X1 U6931 ( .A(\ImageBuffer[24][3] ), .B(\ImageBuffer[25][3] ), .C(
        \ImageBuffer[26][3] ), .D(\ImageBuffer[27][3] ), .S0(n3489), .S1(n3925), .Y(n3831) );
  MX4X1 U6932 ( .A(n3853), .B(n3851), .C(n3852), .D(n3850), .S0(n3933), .S1(
        n3409), .Y(n3854) );
  MX4X1 U6933 ( .A(\ImageBuffer[28][4] ), .B(\ImageBuffer[29][4] ), .C(
        \ImageBuffer[30][4] ), .D(\ImageBuffer[31][4] ), .S0(n3486), .S1(n3924), .Y(n3850) );
  MX4X1 U6934 ( .A(\ImageBuffer[20][4] ), .B(\ImageBuffer[21][4] ), .C(
        \ImageBuffer[22][4] ), .D(\ImageBuffer[23][4] ), .S0(n3486), .S1(n3920), .Y(n3852) );
  MX4X1 U6935 ( .A(\ImageBuffer[24][4] ), .B(\ImageBuffer[25][4] ), .C(
        \ImageBuffer[26][4] ), .D(\ImageBuffer[27][4] ), .S0(n3486), .S1(n3920), .Y(n3851) );
  MX4X1 U6936 ( .A(n3793), .B(n3791), .C(n3792), .D(n3790), .S0(n3933), .S1(
        n3409), .Y(n3794) );
  MX4X1 U6937 ( .A(\ImageBuffer[16][1] ), .B(\ImageBuffer[17][1] ), .C(
        \ImageBuffer[18][1] ), .D(\ImageBuffer[19][1] ), .S0(n3486), .S1(n3932), .Y(n3793) );
  MX4X1 U6938 ( .A(\ImageBuffer[24][1] ), .B(\ImageBuffer[25][1] ), .C(
        \ImageBuffer[26][1] ), .D(\ImageBuffer[27][1] ), .S0(n3486), .S1(n3341), .Y(n3791) );
  MX4X1 U6939 ( .A(\ImageBuffer[28][1] ), .B(\ImageBuffer[29][1] ), .C(
        \ImageBuffer[30][1] ), .D(\ImageBuffer[31][1] ), .S0(n3486), .S1(n3499), .Y(n3790) );
  MX4X1 U6940 ( .A(\ImageBuffer[48][3] ), .B(\ImageBuffer[49][3] ), .C(
        \ImageBuffer[50][3] ), .D(\ImageBuffer[51][3] ), .S0(n3935), .S1(n4303), .Y(n4200) );
  MX4X1 U6941 ( .A(\ImageBuffer[32][3] ), .B(\ImageBuffer[33][3] ), .C(
        \ImageBuffer[34][3] ), .D(\ImageBuffer[35][3] ), .S0(n3935), .S1(n4309), .Y(n4205) );
  MX4X1 U6942 ( .A(\ImageBuffer[28][3] ), .B(\ImageBuffer[29][3] ), .C(
        \ImageBuffer[30][3] ), .D(\ImageBuffer[31][3] ), .S0(n4298), .S1(n4309), .Y(n4207) );
  MX4X1 U6943 ( .A(\ImageBuffer[12][3] ), .B(\ImageBuffer[13][3] ), .C(
        \ImageBuffer[14][3] ), .D(\ImageBuffer[15][3] ), .S0(n4298), .S1(n4310), .Y(n4212) );
  MX4X1 U6944 ( .A(\ImageBuffer[44][3] ), .B(\ImageBuffer[45][3] ), .C(
        \ImageBuffer[46][3] ), .D(\ImageBuffer[47][3] ), .S0(n4298), .S1(n4315), .Y(n4202) );
  MX4X1 U6945 ( .A(\ImageBuffer[8][3] ), .B(\ImageBuffer[9][3] ), .C(
        \ImageBuffer[10][3] ), .D(\ImageBuffer[11][3] ), .S0(n3935), .S1(n4305), .Y(n4213) );
  MX4X1 U6946 ( .A(\ImageBuffer[40][3] ), .B(\ImageBuffer[41][3] ), .C(
        \ImageBuffer[42][3] ), .D(\ImageBuffer[43][3] ), .S0(n3935), .S1(n4307), .Y(n4203) );
  MX4X1 U6947 ( .A(\ImageBuffer[52][3] ), .B(\ImageBuffer[53][3] ), .C(
        \ImageBuffer[54][3] ), .D(\ImageBuffer[55][3] ), .S0(n4298), .S1(n4311), .Y(n4199) );
  MX4X1 U6948 ( .A(\ImageBuffer[4][3] ), .B(\ImageBuffer[5][3] ), .C(
        \ImageBuffer[6][3] ), .D(\ImageBuffer[7][3] ), .S0(n4298), .S1(n4310), 
        .Y(n4214) );
  MX4X1 U6949 ( .A(\ImageBuffer[36][3] ), .B(\ImageBuffer[37][3] ), .C(
        \ImageBuffer[38][3] ), .D(\ImageBuffer[39][3] ), .S0(n4298), .S1(n4313), .Y(n4204) );
  MX4X1 U6950 ( .A(\ImageBuffer[20][7] ), .B(\ImageBuffer[21][7] ), .C(
        \ImageBuffer[22][7] ), .D(\ImageBuffer[23][7] ), .S0(n4119), .S1(n3750), .Y(n4100) );
  MX4X1 U6951 ( .A(\ImageBuffer[4][7] ), .B(\ImageBuffer[5][7] ), .C(
        \ImageBuffer[6][7] ), .D(\ImageBuffer[7][7] ), .S0(n4119), .S1(n3756), 
        .Y(n4105) );
  MX4X1 U6952 ( .A(\ImageBuffer[20][7] ), .B(\ImageBuffer[21][7] ), .C(
        \ImageBuffer[22][7] ), .D(\ImageBuffer[23][7] ), .S0(n3744), .S1(n3757), .Y(n3725) );
  MX4X1 U6953 ( .A(\ImageBuffer[36][7] ), .B(\ImageBuffer[37][7] ), .C(
        \ImageBuffer[38][7] ), .D(\ImageBuffer[39][7] ), .S0(n3744), .S1(n3748), .Y(n3720) );
  MX4X1 U6954 ( .A(\ImageBuffer[4][7] ), .B(\ImageBuffer[5][7] ), .C(
        \ImageBuffer[6][7] ), .D(\ImageBuffer[7][7] ), .S0(n3744), .S1(n3753), 
        .Y(n3730) );
  MX4X1 U6955 ( .A(\ImageBuffer[4][7] ), .B(\ImageBuffer[5][7] ), .C(
        \ImageBuffer[6][7] ), .D(\ImageBuffer[7][7] ), .S0(n3938), .S1(n5123), 
        .Y(n3917) );
  MX4X1 U6956 ( .A(\ImageBuffer[36][7] ), .B(\ImageBuffer[37][7] ), .C(
        \ImageBuffer[38][7] ), .D(\ImageBuffer[39][7] ), .S0(n3938), .S1(n3480), .Y(n3907) );
  MX4X1 U6957 ( .A(\ImageBuffer[20][7] ), .B(\ImageBuffer[21][7] ), .C(
        \ImageBuffer[22][7] ), .D(\ImageBuffer[23][7] ), .S0(n3939), .S1(n4316), .Y(n4289) );
  MX4X1 U6958 ( .A(\ImageBuffer[4][7] ), .B(\ImageBuffer[5][7] ), .C(
        \ImageBuffer[6][7] ), .D(\ImageBuffer[7][7] ), .S0(n3939), .S1(n4311), 
        .Y(n4294) );
  MX4X1 U6959 ( .A(\ImageBuffer[36][7] ), .B(\ImageBuffer[37][7] ), .C(
        \ImageBuffer[38][7] ), .D(\ImageBuffer[39][7] ), .S0(n3939), .S1(n4307), .Y(n4284) );
  MX4X1 U6960 ( .A(\ImageBuffer[0][7] ), .B(\ImageBuffer[1][7] ), .C(
        \ImageBuffer[2][7] ), .D(\ImageBuffer[3][7] ), .S0(n4119), .S1(n3750), 
        .Y(n4106) );
  MX4X1 U6961 ( .A(\ImageBuffer[32][7] ), .B(\ImageBuffer[33][7] ), .C(
        \ImageBuffer[34][7] ), .D(\ImageBuffer[35][7] ), .S0(n3744), .S1(n4128), .Y(n3721) );
  MX4X1 U6962 ( .A(\ImageBuffer[0][7] ), .B(\ImageBuffer[1][7] ), .C(
        \ImageBuffer[2][7] ), .D(\ImageBuffer[3][7] ), .S0(n3744), .S1(n3756), 
        .Y(n3731) );
  MX4X1 U6963 ( .A(\ImageBuffer[0][7] ), .B(\ImageBuffer[1][7] ), .C(
        \ImageBuffer[2][7] ), .D(\ImageBuffer[3][7] ), .S0(n3938), .S1(n3931), 
        .Y(n3918) );
  MX4X1 U6964 ( .A(\ImageBuffer[32][7] ), .B(\ImageBuffer[33][7] ), .C(
        \ImageBuffer[34][7] ), .D(\ImageBuffer[35][7] ), .S0(n3938), .S1(n3930), .Y(n3908) );
  MX4X1 U6965 ( .A(\ImageBuffer[48][7] ), .B(\ImageBuffer[49][7] ), .C(
        \ImageBuffer[50][7] ), .D(\ImageBuffer[51][7] ), .S0(n3939), .S1(n4316), .Y(n4280) );
  MX4X1 U6966 ( .A(\ImageBuffer[0][7] ), .B(\ImageBuffer[1][7] ), .C(
        \ImageBuffer[2][7] ), .D(\ImageBuffer[3][7] ), .S0(n3939), .S1(n4305), 
        .Y(n4295) );
  MX4X1 U6967 ( .A(\ImageBuffer[32][7] ), .B(\ImageBuffer[33][7] ), .C(
        \ImageBuffer[34][7] ), .D(\ImageBuffer[35][7] ), .S0(n3939), .S1(n4304), .Y(n4285) );
  MX4X1 U6968 ( .A(\ImageBuffer[16][7] ), .B(\ImageBuffer[17][7] ), .C(
        \ImageBuffer[18][7] ), .D(\ImageBuffer[19][7] ), .S0(n4119), .S1(n3752), .Y(n4101) );
  MX4X1 U6969 ( .A(\ImageBuffer[24][7] ), .B(\ImageBuffer[25][7] ), .C(
        \ImageBuffer[26][7] ), .D(\ImageBuffer[27][7] ), .S0(n4119), .S1(n3751), .Y(n4099) );
  MX4X1 U6970 ( .A(n3686), .B(n3684), .C(n3685), .D(n3683), .S0(n3734), .S1(
        n3759), .Y(n3687) );
  MX4X1 U6971 ( .A(\ImageBuffer[16][7] ), .B(\ImageBuffer[17][7] ), .C(
        \ImageBuffer[18][7] ), .D(\ImageBuffer[19][7] ), .S0(n3744), .S1(n4122), .Y(n3726) );
  MX4X1 U6972 ( .A(\ImageBuffer[24][7] ), .B(\ImageBuffer[25][7] ), .C(
        \ImageBuffer[26][7] ), .D(\ImageBuffer[27][7] ), .S0(n3744), .S1(n3755), .Y(n3724) );
  MX4X1 U6973 ( .A(\ImageBuffer[28][7] ), .B(\ImageBuffer[29][7] ), .C(
        \ImageBuffer[30][7] ), .D(\ImageBuffer[31][7] ), .S0(n3744), .S1(n4123), .Y(n3723) );
  MX4X1 U6974 ( .A(\ImageBuffer[12][7] ), .B(\ImageBuffer[13][7] ), .C(
        \ImageBuffer[14][7] ), .D(\ImageBuffer[15][7] ), .S0(n4119), .S1(n4132), .Y(n4103) );
  MX4X1 U6975 ( .A(\ImageBuffer[44][7] ), .B(\ImageBuffer[45][7] ), .C(
        \ImageBuffer[46][7] ), .D(\ImageBuffer[47][7] ), .S0(n3744), .S1(n4125), .Y(n3718) );
  MX4X1 U6976 ( .A(\ImageBuffer[12][7] ), .B(\ImageBuffer[13][7] ), .C(
        \ImageBuffer[14][7] ), .D(\ImageBuffer[15][7] ), .S0(n3744), .S1(n5116), .Y(n3728) );
  MX4X1 U6977 ( .A(\ImageBuffer[12][7] ), .B(\ImageBuffer[13][7] ), .C(
        \ImageBuffer[14][7] ), .D(\ImageBuffer[15][7] ), .S0(n3938), .S1(n3920), .Y(n3915) );
  MX4X1 U6978 ( .A(\ImageBuffer[44][7] ), .B(\ImageBuffer[45][7] ), .C(
        \ImageBuffer[46][7] ), .D(\ImageBuffer[47][7] ), .S0(n3938), .S1(n3921), .Y(n3905) );
  MX4X1 U6979 ( .A(\ImageBuffer[12][7] ), .B(\ImageBuffer[13][7] ), .C(
        \ImageBuffer[14][7] ), .D(\ImageBuffer[15][7] ), .S0(n3939), .S1(n4308), .Y(n4292) );
  MX4X1 U6980 ( .A(\ImageBuffer[44][7] ), .B(\ImageBuffer[45][7] ), .C(
        \ImageBuffer[46][7] ), .D(\ImageBuffer[47][7] ), .S0(n3497), .S1(n4316), .Y(n4282) );
  MX4X1 U6981 ( .A(n3716), .B(n3714), .C(n3715), .D(n3713), .S0(n3734), .S1(
        n3759), .Y(n3717) );
  MX4X1 U6982 ( .A(\ImageBuffer[48][7] ), .B(\ImageBuffer[49][7] ), .C(
        \ImageBuffer[50][7] ), .D(\ImageBuffer[51][7] ), .S0(n3744), .S1(n5116), .Y(n3716) );
  MX4X1 U6983 ( .A(\ImageBuffer[56][7] ), .B(\ImageBuffer[57][7] ), .C(
        \ImageBuffer[58][7] ), .D(\ImageBuffer[59][7] ), .S0(n3741), .S1(n3756), .Y(n3714) );
  MX4X1 U6984 ( .A(\ImageBuffer[60][7] ), .B(\ImageBuffer[61][7] ), .C(
        \ImageBuffer[62][7] ), .D(\ImageBuffer[63][7] ), .S0(n4117), .S1(n3757), .Y(n3713) );
  MX4X1 U6985 ( .A(\ImageBuffer[8][7] ), .B(\ImageBuffer[9][7] ), .C(
        \ImageBuffer[10][7] ), .D(\ImageBuffer[11][7] ), .S0(n4119), .S1(n4131), .Y(n4104) );
  MX4X1 U6986 ( .A(\ImageBuffer[40][7] ), .B(\ImageBuffer[41][7] ), .C(
        \ImageBuffer[42][7] ), .D(\ImageBuffer[43][7] ), .S0(n3744), .S1(n4125), .Y(n3719) );
  MX4X1 U6987 ( .A(\ImageBuffer[8][7] ), .B(\ImageBuffer[9][7] ), .C(
        \ImageBuffer[10][7] ), .D(\ImageBuffer[11][7] ), .S0(n3744), .S1(n4127), .Y(n3729) );
  MX4X1 U6988 ( .A(\ImageBuffer[8][7] ), .B(\ImageBuffer[9][7] ), .C(
        \ImageBuffer[10][7] ), .D(\ImageBuffer[11][7] ), .S0(n3938), .S1(n3920), .Y(n3916) );
  MX4X1 U6989 ( .A(\ImageBuffer[40][7] ), .B(\ImageBuffer[41][7] ), .C(
        \ImageBuffer[42][7] ), .D(\ImageBuffer[43][7] ), .S0(n3938), .S1(n3920), .Y(n3906) );
  MX4X1 U6990 ( .A(\ImageBuffer[8][7] ), .B(\ImageBuffer[9][7] ), .C(
        \ImageBuffer[10][7] ), .D(\ImageBuffer[11][7] ), .S0(n3497), .S1(n4307), .Y(n4293) );
  MX4X1 U6991 ( .A(\ImageBuffer[40][7] ), .B(\ImageBuffer[41][7] ), .C(
        \ImageBuffer[42][7] ), .D(\ImageBuffer[43][7] ), .S0(n3939), .S1(n4311), .Y(n4283) );
  MX4X1 U6992 ( .A(\ImageBuffer[32][7] ), .B(\ImageBuffer[33][7] ), .C(
        \ImageBuffer[34][7] ), .D(\ImageBuffer[35][7] ), .S0(n4119), .S1(n4132), .Y(n4096) );
  MX4X1 U6993 ( .A(\ImageBuffer[40][7] ), .B(\ImageBuffer[41][7] ), .C(
        \ImageBuffer[42][7] ), .D(\ImageBuffer[43][7] ), .S0(n4119), .S1(n3753), .Y(n4094) );
  MX4X1 U6994 ( .A(\ImageBuffer[44][7] ), .B(\ImageBuffer[45][7] ), .C(
        \ImageBuffer[46][7] ), .D(\ImageBuffer[47][7] ), .S0(n4119), .S1(n4130), .Y(n4093) );
  MX4X1 U6995 ( .A(\ImageBuffer[28][7] ), .B(\ImageBuffer[29][7] ), .C(
        \ImageBuffer[30][7] ), .D(\ImageBuffer[31][7] ), .S0(n3938), .S1(n3920), .Y(n3910) );
  MX4X1 U6996 ( .A(\ImageBuffer[20][7] ), .B(\ImageBuffer[21][7] ), .C(
        \ImageBuffer[22][7] ), .D(\ImageBuffer[23][7] ), .S0(n3938), .S1(n3930), .Y(n3912) );
  INVX3 U6997 ( .A(reset), .Y(n8602) );
  ADDHXL U6998 ( .A(n8621), .B(n8622), .CO(\add_122/carry[2] ), .S(N2545) );
  ADDHXL U6999 ( .A(IROM_A[3]), .B(\add_122/carry[3] ), .CO(\add_122/carry[4] ), .S(N2547) );
  ADDHXL U7000 ( .A(n8620), .B(\add_122/carry[2] ), .CO(\add_122/carry[3] ), 
        .S(N2546) );
  ADDHXL U7001 ( .A(IROM_A[4]), .B(\add_122/carry[4] ), .CO(\add_122/carry[5] ), .S(N2548) );
  MX4X1 U7002 ( .A(n4655), .B(n4653), .C(n4654), .D(n4652), .S0(N2520), .S1(
        n4819), .Y(n4656) );
  MX4X1 U7003 ( .A(n4675), .B(n4673), .C(n4674), .D(n4672), .S0(n4820), .S1(
        n4818), .Y(n4676) );
  MX4X1 U7004 ( .A(n4695), .B(n4693), .C(n4694), .D(n4692), .S0(n4820), .S1(
        n4818), .Y(n4696) );
  MX4X1 U7005 ( .A(n4715), .B(n4713), .C(n4714), .D(n4712), .S0(n4820), .S1(
        n4818), .Y(n4716) );
  MX4X1 U7006 ( .A(n4735), .B(n4733), .C(n4734), .D(n4732), .S0(n4820), .S1(
        n4818), .Y(n4736) );
  MX4X1 U7007 ( .A(n4755), .B(n4753), .C(n4754), .D(n4752), .S0(n4821), .S1(
        n4819), .Y(n4756) );
  MX4X1 U7008 ( .A(n4775), .B(n4773), .C(n4774), .D(n4772), .S0(n4821), .S1(
        n4819), .Y(n4776) );
  MX4X1 U7009 ( .A(n4795), .B(n4793), .C(n4794), .D(n4792), .S0(n4821), .S1(
        n4819), .Y(n4796) );
  MX4X1 U7010 ( .A(n4661), .B(n4651), .C(n4656), .D(n4646), .S0(N2522), .S1(
        N2521), .Y(N13071) );
  MX4X1 U7011 ( .A(n4650), .B(n4648), .C(n4649), .D(n4647), .S0(N2520), .S1(
        n4819), .Y(n4651) );
  MX4X1 U7012 ( .A(n4645), .B(n4643), .C(n4644), .D(n4642), .S0(n5104), .S1(
        n4818), .Y(n4646) );
  MX4X1 U7013 ( .A(n4660), .B(n4658), .C(n4659), .D(n4657), .S0(n5104), .S1(
        n4819), .Y(n4661) );
  MX4X1 U7014 ( .A(n4681), .B(n4671), .C(n4676), .D(n4666), .S0(N2522), .S1(
        N2521), .Y(N13070) );
  MX4X1 U7015 ( .A(n4680), .B(n4678), .C(n4679), .D(n4677), .S0(n4820), .S1(
        n4818), .Y(n4681) );
  MX4X1 U7016 ( .A(n4670), .B(n4668), .C(n4669), .D(n4667), .S0(n5104), .S1(
        n4818), .Y(n4671) );
  MX4X1 U7017 ( .A(n4665), .B(n4663), .C(n4664), .D(n4662), .S0(N2520), .S1(
        n4818), .Y(n4666) );
  MX4X1 U7018 ( .A(n4701), .B(n4691), .C(n4696), .D(n4686), .S0(N2522), .S1(
        N2521), .Y(N13069) );
  MX4X1 U7019 ( .A(n4700), .B(n4698), .C(n4699), .D(n4697), .S0(n4820), .S1(
        n4818), .Y(n4701) );
  MX4X1 U7020 ( .A(n4690), .B(n4688), .C(n4689), .D(n4687), .S0(n4820), .S1(
        n4818), .Y(n4691) );
  MX4X1 U7021 ( .A(n4685), .B(n4683), .C(n4684), .D(n4682), .S0(n4820), .S1(
        n4818), .Y(n4686) );
  MX4X1 U7022 ( .A(n4721), .B(n4711), .C(n4716), .D(n4706), .S0(N2522), .S1(
        N2521), .Y(N13068) );
  MX4X1 U7023 ( .A(n4720), .B(n4718), .C(n4719), .D(n4717), .S0(n4820), .S1(
        n4818), .Y(n4721) );
  MX4X1 U7024 ( .A(n4710), .B(n4708), .C(n4709), .D(n4707), .S0(n4820), .S1(
        n4818), .Y(n4711) );
  MX4X1 U7025 ( .A(n4705), .B(n4703), .C(n4704), .D(n4702), .S0(n4820), .S1(
        n4818), .Y(n4706) );
  MX4X1 U7026 ( .A(n4741), .B(n4731), .C(n4736), .D(n4726), .S0(N2522), .S1(
        N2521), .Y(N13067) );
  MX4X1 U7027 ( .A(n4740), .B(n4738), .C(n4739), .D(n4737), .S0(n4821), .S1(
        n4819), .Y(n4741) );
  MX4X1 U7028 ( .A(n4730), .B(n4728), .C(n4729), .D(n4727), .S0(n4820), .S1(
        n4818), .Y(n4731) );
  MX4X1 U7029 ( .A(n4725), .B(n4723), .C(n4724), .D(n4722), .S0(n4820), .S1(
        n4818), .Y(n4726) );
  MX4X1 U7030 ( .A(n4761), .B(n4751), .C(n4756), .D(n4746), .S0(N2522), .S1(
        N2521), .Y(N13066) );
  MX4X1 U7031 ( .A(n4760), .B(n4758), .C(n4759), .D(n4757), .S0(n4821), .S1(
        n4819), .Y(n4761) );
  MX4X1 U7032 ( .A(n4750), .B(n4748), .C(n4749), .D(n4747), .S0(n4821), .S1(
        n4819), .Y(n4751) );
  MX4X1 U7033 ( .A(n4745), .B(n4743), .C(n4744), .D(n4742), .S0(n4821), .S1(
        n4819), .Y(n4746) );
  MX4X1 U7034 ( .A(n4781), .B(n4771), .C(n4776), .D(n4766), .S0(N2522), .S1(
        N2521), .Y(N13065) );
  MX4X1 U7035 ( .A(n4780), .B(n4778), .C(n4779), .D(n4777), .S0(n4821), .S1(
        n4819), .Y(n4781) );
  MX4X1 U7036 ( .A(n4770), .B(n4768), .C(n4769), .D(n4767), .S0(n4821), .S1(
        n4819), .Y(n4771) );
  MX4X1 U7037 ( .A(n4765), .B(n4763), .C(n4764), .D(n4762), .S0(n4821), .S1(
        n4819), .Y(n4766) );
  MX4X1 U7038 ( .A(n4801), .B(n4791), .C(n4796), .D(n4786), .S0(N2522), .S1(
        N2521), .Y(N13064) );
  MX4X1 U7039 ( .A(n4800), .B(n4798), .C(n4799), .D(n4797), .S0(n4821), .S1(
        n4819), .Y(n4801) );
  MX4X1 U7040 ( .A(n4790), .B(n4788), .C(n4789), .D(n4787), .S0(n4821), .S1(
        n4819), .Y(n4791) );
  MX4X1 U7041 ( .A(n4785), .B(n4783), .C(n4784), .D(n4782), .S0(n4821), .S1(
        n4819), .Y(n4786) );
  CLKBUFX3 U7042 ( .A(N2518), .Y(n5105) );
  CLKBUFX3 U7043 ( .A(N2520), .Y(n5104) );
  ADDHXL U7044 ( .A(N2521), .B(\add_134/carry[4] ), .CO(\add_134/carry[5] ), 
        .S(N2571) );
  MX4X2 U7045 ( .A(n3763), .B(n3761), .C(n3762), .D(n3760), .S0(n3934), .S1(
        n3409), .Y(n3764) );
  MX4X2 U7046 ( .A(n3768), .B(n3766), .C(n3767), .D(n3765), .S0(n3934), .S1(
        n3409), .Y(n3769) );
  MX4X2 U7047 ( .A(n3803), .B(n3801), .C(n3802), .D(n3800), .S0(n3933), .S1(
        N2489), .Y(n3804) );
  MX4X2 U7048 ( .A(n3813), .B(n3811), .C(n3812), .D(n3810), .S0(n3933), .S1(
        N2489), .Y(n3814) );
  MX4X2 U7049 ( .A(n3819), .B(n3809), .C(n3814), .D(n3804), .S0(N2492), .S1(
        N2491), .Y(N2763) );
  MX4X1 U7050 ( .A(n3859), .B(n3849), .C(n3854), .D(n3844), .S0(N2492), .S1(
        N2491), .Y(N2761) );
  MX4XL U7051 ( .A(n3919), .B(n3909), .C(n3914), .D(n3904), .S0(N2492), .S1(
        N2491), .Y(N2758) );
  MX4X1 U7052 ( .A(n3879), .B(n3869), .C(n3874), .D(n3864), .S0(N2492), .S1(
        N2491), .Y(N2760) );
  MX4X2 U7053 ( .A(n4140), .B(n4138), .C(n4139), .D(n4137), .S0(n5108), .S1(
        n3487), .Y(n4141) );
  MX4X2 U7054 ( .A(n4150), .B(n4148), .C(n4149), .D(n4147), .S0(n3493), .S1(
        n3487), .Y(n4151) );
  MX4X2 U7055 ( .A(n4155), .B(n4153), .C(n4154), .D(n4152), .S0(n3493), .S1(
        n3487), .Y(n4156) );
  MX4X2 U7056 ( .A(n4176), .B(n4166), .C(n4171), .D(n4161), .S0(N2504), .S1(
        N2503), .Y(N2772) );
  MX4X2 U7057 ( .A(n4180), .B(n4178), .C(n4179), .D(n4177), .S0(n3493), .S1(
        n3487), .Y(n4181) );
  MX4X2 U7058 ( .A(n4185), .B(n4183), .C(n4184), .D(n4182), .S0(n5108), .S1(
        n3487), .Y(n4186) );
  MX4X2 U7059 ( .A(n4190), .B(n4188), .C(n4189), .D(n4187), .S0(n5108), .S1(
        n3487), .Y(n4191) );
  MX4X2 U7060 ( .A(n4195), .B(n4193), .C(n4194), .D(n4192), .S0(n5108), .S1(
        n3487), .Y(n4196) );
  MX4X2 U7061 ( .A(n4236), .B(n4226), .C(n4231), .D(n4221), .S0(N2504), .S1(
        N2503), .Y(N2769) );
  MX4X2 U7062 ( .A(n4256), .B(n4246), .C(n4251), .D(n4241), .S0(N2504), .S1(
        N2503), .Y(N2768) );
  MX4X2 U7063 ( .A(n4276), .B(n4266), .C(n4271), .D(n4261), .S0(N2504), .S1(
        N2503), .Y(N2767) );
  MX4X2 U7064 ( .A(n4296), .B(n4286), .C(n4291), .D(n4281), .S0(N2504), .S1(
        N2503), .Y(N2766) );
  MX4X4 U7065 ( .A(n4156), .B(n4146), .C(n4151), .D(n4141), .S0(N2504), .S1(
        N2503), .Y(N2773) );
  MX4XL U7066 ( .A(n4210), .B(n4208), .C(n4209), .D(n4207), .S0(n5108), .S1(
        n3487), .Y(n4211) );
  MX4XL U7067 ( .A(n4200), .B(n4198), .C(n4199), .D(n4197), .S0(n5108), .S1(
        n3487), .Y(n4201) );
  MX4XL U7068 ( .A(n4215), .B(n4213), .C(n4214), .D(n4212), .S0(N2502), .S1(
        n3487), .Y(n4216) );
  MX4XL U7069 ( .A(n4205), .B(n4203), .C(n4204), .D(n4202), .S0(n5108), .S1(
        n3487), .Y(n4206) );
  MX4X1 U7070 ( .A(n4338), .B(n4328), .C(n4333), .D(n4323), .S0(N2510), .S1(
        N2509), .Y(N2749) );
  MX4X1 U7071 ( .A(n4398), .B(n4388), .C(n4393), .D(n4383), .S0(N2510), .S1(
        N2509), .Y(N2746) );
  MX4X1 U7072 ( .A(n4518), .B(n4508), .C(n4513), .D(n4503), .S0(N2516), .S1(
        N2515), .Y(N2756) );
  OAI211X1 U7073 ( .A0(n5371), .A1(n5079), .B0(n5370), .C0(n5380), .Y(n5372)
         );
  CLKINVX1 U7074 ( .A(n5319), .Y(n5340) );
  NOR3BX1 U7075 ( .AN(n5334), .B(n5333), .C(n5318), .Y(n5319) );
  CLKBUFX3 U7076 ( .A(n5837), .Y(n4925) );
  CLKINVX1 U7077 ( .A(n5348), .Y(n5369) );
  NOR3BX1 U7078 ( .AN(n5363), .B(n5362), .C(n5347), .Y(n5348) );
  AND2X2 U7079 ( .A(n5253), .B(n5262), .Y(n5259) );
  CLKINVX1 U7080 ( .A(n5256), .Y(n5279) );
  AND2X2 U7081 ( .A(n5283), .B(n5293), .Y(n5290) );
  NAND2BX1 U7082 ( .AN(N2771), .B(n4872), .Y(n5293) );
  CLKINVX1 U7083 ( .A(n5227), .Y(n5249) );
  INVX1 U7084 ( .A(N2771), .Y(n6787) );
  OAI211XL U7085 ( .A0(n5077), .A1(n5382), .B0(n5381), .C0(n5380), .Y(n5384)
         );
  AND2X2 U7086 ( .A(n5373), .B(n5383), .Y(n5380) );
  INVX12 U7087 ( .A(n4945), .Y(N2538) );
  OAI21XL U7088 ( .A0(n5978), .A1(n5979), .B0(n5980), .Y(n8153) );
  NAND2X2 U7089 ( .A(n5043), .B(n4942), .Y(n5979) );
  NAND3BX2 U7090 ( .AN(n5205), .B(n5204), .C(n5203), .Y(n5209) );
  OAI31X1 U7091 ( .A0(n5246), .A1(n5245), .A2(n5244), .B0(n5243), .Y(N2701) );
  AOI31X2 U7092 ( .A0(n5388), .A1(n5373), .A2(n5372), .B0(n5385), .Y(n5375) );
  AOI31X2 U7093 ( .A0(n5398), .A1(n5378), .A2(n5394), .B0(n5397), .Y(n5379) );
  NAND2X6 U7094 ( .A(n8073), .B(n8074), .Y(n8063) );
  CLKINVX1 U7095 ( .A(n5287), .Y(n5311) );
  NOR3BX1 U7096 ( .AN(n5302), .B(n5301), .C(n5286), .Y(n5287) );
  NAND2X2 U7097 ( .A(n7410), .B(n3557), .Y(n7323) );
  NOR4BXL U7098 ( .AN(n8056), .B(n3476), .C(n3477), .D(n3475), .Y(n8060) );
  OAI32X4 U7099 ( .A0(n7739), .A1(n5057), .A2(n7740), .B0(n3352), .B1(n7746), 
        .Y(n7745) );
  OAI32X4 U7100 ( .A0(n7766), .A1(n7192), .A2(n7762), .B0(n5067), .B1(n3368), 
        .Y(n7765) );
  OAI32X4 U7101 ( .A0(n7940), .A1(n5059), .A2(n7941), .B0(n3351), .B1(n7948), 
        .Y(n7947) );
  NAND2XL U7102 ( .A(n7713), .B(n3557), .Y(n7626) );
  OAI32X4 U7103 ( .A0(n7796), .A1(n5057), .A2(n7797), .B0(n3351), .B1(n7803), 
        .Y(n7802) );
  OAI32X4 U7104 ( .A0(n7800), .A1(n7192), .A2(n7796), .B0(n5070), .B1(n3368), 
        .Y(n7799) );
  NAND3X2 U7105 ( .A(n7515), .B(n7717), .C(n5128), .Y(n7833) );
  OAI32X4 U7106 ( .A0(n7215), .A1(n7192), .A2(n7211), .B0(n7193), .B1(n5065), 
        .Y(n7214) );
  OAI32X4 U7107 ( .A0(n7983), .A1(n7192), .A2(n7978), .B0(n3560), .B1(n7928), 
        .Y(n7982) );
  OAI32X4 U7108 ( .A0(n7245), .A1(n7192), .A2(n7241), .B0(n7193), .B1(n5067), 
        .Y(n7244) );
  OAI32X4 U7109 ( .A0(n8006), .A1(n5053), .A2(n8002), .B0(n5070), .B1(n7931), 
        .Y(n8007) );
  OAI32X4 U7110 ( .A0(n8006), .A1(n7192), .A2(n8002), .B0(n5070), .B1(n7928), 
        .Y(n8005) );
  NAND2X2 U7111 ( .A(n8025), .B(n3557), .Y(n7928) );
  OAI33X4 U7112 ( .A0(n7322), .A1(n7192), .A2(n7318), .B0(n7323), .B1(n7324), 
        .B2(n5052), .Y(n7321) );
  OAI32X4 U7113 ( .A0(n7419), .A1(n5055), .A2(n7420), .B0(n3352), .B1(n7427), 
        .Y(n7428) );
  OAI33X4 U7114 ( .A0(n7423), .A1(n7192), .A2(n7419), .B0(n3367), .B1(n7424), 
        .B2(n5052), .Y(n7422) );
  OAI32X4 U7115 ( .A0(n7521), .A1(n5055), .A2(n7522), .B0(n3352), .B1(n7530), 
        .Y(n7531) );
  OAI33X4 U7116 ( .A0(n7525), .A1(n5053), .A2(n7521), .B0(n7529), .B1(n7527), 
        .B2(n5052), .Y(n7528) );
  OAI33X4 U7117 ( .A0(n7350), .A1(n7192), .A2(n7346), .B0(n7323), .B1(n7351), 
        .B2(n3561), .Y(n7349) );
  OAI32X4 U7118 ( .A0(n7446), .A1(n5055), .A2(n7447), .B0(n3351), .B1(n7453), 
        .Y(n7454) );
  OAI33X4 U7119 ( .A0(n7450), .A1(n7192), .A2(n7446), .B0(n3367), .B1(n7451), 
        .B2(n3561), .Y(n7449) );
  OAI32X4 U7120 ( .A0(n7549), .A1(n5056), .A2(n7550), .B0(n3351), .B1(n7556), 
        .Y(n7557) );
  OAI32X4 U7121 ( .A0(n7621), .A1(n5057), .A2(n7622), .B0(n3352), .B1(n7630), 
        .Y(n7631) );
  OAI33X4 U7122 ( .A0(n7826), .A1(n7192), .A2(n7822), .B0(n3369), .B1(n7827), 
        .B2(n3548), .Y(n7825) );
  OAI32X4 U7123 ( .A0(n7583), .A1(n5056), .A2(n7584), .B0(n3351), .B1(n7590), 
        .Y(n7591) );
  OAI32X4 U7124 ( .A0(n7649), .A1(n5056), .A2(n7650), .B0(n3351), .B1(n7656), 
        .Y(n7657) );
  OAI33X4 U7125 ( .A0(n7853), .A1(n7192), .A2(n7849), .B0(n3369), .B1(n7854), 
        .B2(n5066), .Y(n7852) );
  OAI33X4 U7126 ( .A0(n7272), .A1(n7192), .A2(n7268), .B0(n5069), .B1(n7273), 
        .B2(n7193), .Y(n7271) );
  OAI32X4 U7127 ( .A0(n7683), .A1(n5057), .A2(n7684), .B0(n3351), .B1(n7690), 
        .Y(n7691) );
  OAI32X4 U7128 ( .A0(n7883), .A1(n5057), .A2(n7884), .B0(n3352), .B1(n7890), 
        .Y(n7891) );
  OAI33X4 U7129 ( .A0(n7887), .A1(n7192), .A2(n7883), .B0(n3369), .B1(n7888), 
        .B2(n5069), .Y(n7886) );
  OAI33X4 U7130 ( .A0(n7300), .A1(n7192), .A2(n7296), .B0(n5071), .B1(n7301), 
        .B2(n7193), .Y(n7299) );
  OAI32X4 U7131 ( .A0(n7723), .A1(n5057), .A2(n7724), .B0(n3351), .B1(n7731), 
        .Y(n7732) );
  OAI32X4 U7132 ( .A0(n7750), .A1(n5057), .A2(n7751), .B0(n3352), .B1(n7757), 
        .Y(n7758) );
  OAI32X4 U7133 ( .A0(n8016), .A1(n5059), .A2(n8017), .B0(n3352), .B1(n8027), 
        .Y(n8032) );
  OAI33X4 U7134 ( .A0(n8023), .A1(n7192), .A2(n8016), .B0(n7928), .B1(n8024), 
        .B2(n3558), .Y(n8022) );
  OAI32X4 U7135 ( .A0(n7784), .A1(n5058), .A2(n7785), .B0(n3352), .B1(n7791), 
        .Y(n7792) );
  OAI33X4 U7136 ( .A0(n7788), .A1(n7192), .A2(n7784), .B0(n3368), .B1(n7789), 
        .B2(n3562), .Y(n7787) );
  OAI33X4 U7137 ( .A0(n7927), .A1(n7192), .A2(n7920), .B0(n7928), .B1(n7929), 
        .B2(n3548), .Y(n7926) );
  OAI31X2 U7138 ( .A0(n5217), .A1(n5216), .A2(n5215), .B0(n5214), .Y(N2697) );
  AOI31X4 U7139 ( .A0(N2703), .A1(N2701), .A2(N2702), .B0(n8065), .Y(n8073) );
  AOI211X2 U7140 ( .A0(n5213), .A1(n5212), .B0(n5211), .C0(n5210), .Y(n5215)
         );
  OAI221X4 U7141 ( .A0(n7515), .A1(n8076), .B0(n7310), .B1(n8077), .C0(n8081), 
        .Y(N2509) );
  AOI2BB2XL U7142 ( .B0(n8065), .B1(n5125), .A0N(n7307), .A1N(n3523), .Y(n8067) );
  OAI221X4 U7143 ( .A0(n7515), .A1(n3348), .B0(n7310), .B1(n8063), .C0(n8067), 
        .Y(N2515) );
  OAI221X4 U7144 ( .A0(n7717), .A1(n3348), .B0(n7311), .B1(n8063), .C0(n8064), 
        .Y(N2516) );
  AOI31X4 U7145 ( .A0(N2675), .A1(N2673), .A2(N2674), .B0(n8079), .Y(n8086) );
  NOR3BX2 U7146 ( .AN(n5180), .B(n5179), .C(n5164), .Y(n5165) );
  OAI221X4 U7147 ( .A0(n7717), .A1(n8076), .B0(n7311), .B1(n8077), .C0(n8078), 
        .Y(N2510) );
  NOR3BX2 U7148 ( .AN(n5212), .B(n5211), .C(n5196), .Y(n5197) );
  CLKXOR2X8 U7149 ( .A(n4947), .B(\add_80/carry[5] ), .Y(N2504) );
  XNOR2X1 U7150 ( .A(n4947), .B(\sub_157_S2_aco/carry[5] ), .Y(N2615) );
  XNOR2X1 U7151 ( .A(\sub_157_S2_aco/carry[4] ), .B(n5125), .Y(N2614) );
  OR2X1 U7152 ( .A(n3371), .B(n5127), .Y(\sub_157_S2_aco/carry[4] ) );
  XNOR2X1 U7153 ( .A(n5127), .B(n3371), .Y(N2613) );
  XNOR2X1 U7154 ( .A(n4947), .B(\sub_168_aco/carry[5] ), .Y(N2635) );
  XNOR2X1 U7155 ( .A(\sub_168_aco/carry[4] ), .B(n5125), .Y(N2634) );
  OR2X1 U7156 ( .A(n5127), .B(\sub_168_aco/carry[3] ), .Y(
        \sub_168_aco/carry[4] ) );
  XNOR2X1 U7157 ( .A(\sub_168_aco/carry[3] ), .B(n5127), .Y(N2633) );
  OR2X1 U7158 ( .A(N2495), .B(\sub_168_aco/carry[2] ), .Y(
        \sub_168_aco/carry[3] ) );
  OR2X1 U7159 ( .A(n4134), .B(\sub_168_aco/carry[1] ), .Y(
        \sub_168_aco/carry[2] ) );
  XNOR2X1 U7160 ( .A(\sub_168_aco/carry[1] ), .B(n4123), .Y(N2631) );
  XOR2X1 U7161 ( .A(n4947), .B(\add_162_S2_aco/carry[5] ), .Y(N2625) );
  AND2X1 U7162 ( .A(\add_162_S2_aco/carry[4] ), .B(n5125), .Y(
        \add_162_S2_aco/carry[5] ) );
  AND2X1 U7163 ( .A(n5127), .B(N2617), .Y(\add_162_S2_aco/carry[4] ) );
  XOR2X1 U7164 ( .A(N2617), .B(n5127), .Y(N2623) );
  OR2X1 U7165 ( .A(n7295), .B(n5118), .Y(\sub_168_aco/carry[1] ) );
  XNOR2X1 U7166 ( .A(n5118), .B(n7295), .Y(N2630) );
  XOR2X1 U7167 ( .A(\add_134/carry[5] ), .B(N2522), .Y(N2572) );
  NAND2BX1 U7168 ( .AN(n4869), .B(n4863), .Y(n5149) );
  NAND2X1 U7169 ( .A(n4868), .B(n5219), .Y(n5136) );
  NAND2X1 U7170 ( .A(n4871), .B(n5156), .Y(n5145) );
  NAND2BX1 U7171 ( .AN(N2779), .B(n4872), .Y(n5131) );
  NAND2BX1 U7172 ( .AN(n4872), .B(N2779), .Y(n5140) );
  NOR2X1 U7173 ( .A(n5156), .B(N2762), .Y(n5142) );
  OAI2BB1X1 U7174 ( .A0N(n5222), .A1N(n4866), .B0(n4873), .Y(n5139) );
  OAI211X1 U7175 ( .A0(n4866), .A1(n5222), .B0(n5139), .C0(n5138), .Y(n5141)
         );
  NAND3BX1 U7176 ( .AN(n5142), .B(n5141), .C(n5140), .Y(n5146) );
  NAND2X1 U7177 ( .A(n5096), .B(n5187), .Y(n5166) );
  NOR2BX1 U7178 ( .AN(n5091), .B(n4864), .Y(n5162) );
  NAND2X1 U7179 ( .A(n5101), .B(n5188), .Y(n5182) );
  OAI2BB1X1 U7180 ( .A0N(n5170), .A1N(n4866), .B0(n5077), .Y(n5169) );
  OAI211X1 U7181 ( .A0(n4866), .A1(n5170), .B0(n5169), .C0(n5168), .Y(n5172)
         );
  NAND3BX1 U7182 ( .AN(n5173), .B(n5172), .C(n5171), .Y(n5177) );
  CLKINVX6 U7183 ( .A(n5165), .Y(n5189) );
  NAND2BX1 U7184 ( .AN(N2768), .B(n4863), .Y(n5212) );
  NAND2BX1 U7185 ( .AN(n5216), .B(n5198), .Y(n5211) );
  NAND2BX1 U7186 ( .AN(N2779), .B(N2771), .Y(n5193) );
  NAND2BX1 U7187 ( .AN(N2771), .B(N2779), .Y(n5203) );
  AOI31X1 U7188 ( .A0(n5208), .A1(n5193), .A2(n5192), .B0(n5205), .Y(n5195) );
  NOR2BX1 U7189 ( .AN(N2769), .B(n4864), .Y(n5194) );
  NOR2BX1 U7190 ( .AN(n4864), .B(N2769), .Y(n5206) );
  NAND2X1 U7191 ( .A(N2766), .B(n5157), .Y(n5214) );
  NOR2BX1 U7192 ( .AN(N2781), .B(N2773), .Y(n5202) );
  OAI2BB1X1 U7193 ( .A0N(n5202), .A1N(n4866), .B0(N2772), .Y(n5201) );
  NOR2X1 U7194 ( .A(n5248), .B(n4862), .Y(n5245) );
  NAND2X1 U7195 ( .A(n4862), .B(n5248), .Y(n5228) );
  NAND2BX1 U7196 ( .AN(n4872), .B(N2779), .Y(n5224) );
  NAND2BX1 U7197 ( .AN(N2779), .B(n4872), .Y(n5233) );
  AND2X1 U7198 ( .A(n5224), .B(n5233), .Y(n5230) );
  AOI31X1 U7199 ( .A0(n5237), .A1(n5224), .A2(n5223), .B0(n5235), .Y(n5225) );
  NOR2X1 U7200 ( .A(n5143), .B(n5132), .Y(n5236) );
  AOI211X1 U7201 ( .A0(n5225), .A1(n5236), .B0(n5143), .C0(n5239), .Y(n5226)
         );
  NAND2X1 U7202 ( .A(n4861), .B(n5250), .Y(n5243) );
  AOI31X1 U7203 ( .A0(n5249), .A1(n5228), .A2(n5243), .B0(n5246), .Y(n5229) );
  OAI2BB1X1 U7204 ( .A0N(n5232), .A1N(n4873), .B0(n4866), .Y(n5231) );
  OAI211X1 U7205 ( .A0(n4873), .A1(n5232), .B0(n5231), .C0(n5230), .Y(n5234)
         );
  NAND3BX1 U7206 ( .AN(n5235), .B(n5234), .C(n5233), .Y(n5238) );
  AOI31X1 U7207 ( .A0(n5238), .A1(n5237), .A2(n5236), .B0(n5132), .Y(n5242) );
  AOI211X1 U7208 ( .A0(n5242), .A1(n5241), .B0(n5240), .C0(n5239), .Y(n5244)
         );
  NOR2X1 U7209 ( .A(n5278), .B(n5096), .Y(n5274) );
  NAND2X1 U7210 ( .A(n5096), .B(n5278), .Y(n5257) );
  AO21X1 U7211 ( .A0(n5276), .A1(n5353), .B0(n5077), .Y(n5251) );
  OAI211X1 U7212 ( .A0(n5353), .A1(n5276), .B0(n5251), .C0(n5259), .Y(n5252)
         );
  NOR2X1 U7213 ( .A(n5357), .B(n3492), .Y(n5265) );
  NAND2X1 U7214 ( .A(n5101), .B(n5250), .Y(n5272) );
  AOI31X1 U7215 ( .A0(n5279), .A1(n5257), .A2(n5272), .B0(n5275), .Y(n5258) );
  NOR2X1 U7216 ( .A(n5278), .B(N2767), .Y(n5306) );
  NAND2X1 U7217 ( .A(N2767), .B(n5278), .Y(n5288) );
  NAND2X1 U7218 ( .A(N2770), .B(n5309), .Y(n5298) );
  NAND2BX1 U7219 ( .AN(n4872), .B(N2771), .Y(n5283) );
  NOR2BX1 U7220 ( .AN(N2773), .B(N2765), .Y(n5281) );
  AO21X1 U7221 ( .A0(n5308), .A1(n5281), .B0(N2772), .Y(n5280) );
  OAI211X1 U7222 ( .A0(n5281), .A1(n5308), .B0(n5280), .C0(n5290), .Y(n5282)
         );
  NOR2X1 U7223 ( .A(n5309), .B(N2770), .Y(n5295) );
  NOR2BX1 U7224 ( .AN(N2769), .B(n4870), .Y(n5284) );
  NOR2BX1 U7225 ( .AN(n4870), .B(N2769), .Y(n5296) );
  NOR2BX1 U7226 ( .AN(N2768), .B(n4869), .Y(n5300) );
  NAND2X1 U7227 ( .A(N2766), .B(n5310), .Y(n5304) );
  NOR2BX1 U7228 ( .AN(N2765), .B(N2773), .Y(n5292) );
  OAI2BB1X1 U7229 ( .A0N(n5292), .A1N(n4873), .B0(N2772), .Y(n5291) );
  OAI211X1 U7230 ( .A0(n4873), .A1(n5292), .B0(n5291), .C0(n5290), .Y(n5294)
         );
  AOI31X1 U7231 ( .A0(n5299), .A1(n5298), .A2(n5297), .B0(n5296), .Y(n5303) );
  AOI211X1 U7232 ( .A0(n5303), .A1(n5302), .B0(n5301), .C0(n5300), .Y(n5305)
         );
  NOR2X1 U7233 ( .A(n5097), .B(n4862), .Y(n5338) );
  NAND2X1 U7234 ( .A(n4862), .B(n5097), .Y(n5320) );
  NAND2BX1 U7235 ( .AN(n3944), .B(N2779), .Y(n5315) );
  NOR2BX1 U7236 ( .AN(N2781), .B(n5074), .Y(n5313) );
  NAND2BX1 U7237 ( .AN(N2779), .B(n3944), .Y(n5325) );
  OAI211X1 U7238 ( .A0(n5313), .A1(n5078), .B0(n5312), .C0(n5322), .Y(n5314)
         );
  AOI31X1 U7239 ( .A0(n5330), .A1(n5315), .A2(n5314), .B0(n5327), .Y(n5317) );
  AOI211X1 U7240 ( .A0(n5317), .A1(n5329), .B0(n5316), .C0(n5332), .Y(n5318)
         );
  NAND2X1 U7241 ( .A(n4861), .B(n5102), .Y(n5336) );
  AOI31X1 U7242 ( .A0(n5340), .A1(n5320), .A2(n5336), .B0(n5339), .Y(n5321) );
  AOI211X1 U7243 ( .A0(n5335), .A1(n5334), .B0(n5333), .C0(n5332), .Y(n5337)
         );
  NAND2BX1 U7244 ( .AN(n4869), .B(n5093), .Y(n5363) );
  NOR2X1 U7245 ( .A(n5097), .B(n4868), .Y(n5367) );
  NAND2X1 U7246 ( .A(n4868), .B(n5098), .Y(n5349) );
  NAND2X1 U7247 ( .A(n4871), .B(n5086), .Y(n5359) );
  NAND2BX1 U7248 ( .AN(n3944), .B(n4872), .Y(n5344) );
  NOR2BX1 U7249 ( .AN(N2765), .B(n5074), .Y(n5342) );
  NAND2BX1 U7250 ( .AN(n4872), .B(n3944), .Y(n5354) );
  NOR2X1 U7251 ( .A(n5087), .B(n4871), .Y(n5356) );
  AOI31X1 U7252 ( .A0(n5359), .A1(n5344), .A2(n5343), .B0(n5356), .Y(n5346) );
  NOR2BX1 U7253 ( .AN(n4869), .B(n5093), .Y(n5361) );
  AOI211X1 U7254 ( .A0(n5346), .A1(n5358), .B0(n3492), .C0(n5361), .Y(n5347)
         );
  NAND2X1 U7255 ( .A(n4867), .B(n5102), .Y(n5365) );
  NOR2X1 U7256 ( .A(n5102), .B(n4867), .Y(n5368) );
  AOI31X1 U7257 ( .A0(n5369), .A1(n5349), .A2(n5365), .B0(n5368), .Y(n5350) );
  AOI211X1 U7258 ( .A0(n5364), .A1(n5363), .B0(n5362), .C0(n5361), .Y(n5366)
         );
  NAND2X1 U7259 ( .A(N2770), .B(n5087), .Y(n5388) );
  NOR2X1 U7260 ( .A(n5086), .B(N2770), .Y(n5385) );
  NOR2X1 U7261 ( .A(n5374), .B(n5386), .Y(n5387) );
  NOR2BX1 U7262 ( .AN(n5074), .B(N2773), .Y(n5382) );
  OAI2BB1X1 U7263 ( .A0N(n5382), .A1N(n5077), .B0(N2772), .Y(n5381) );
  NAND3BX1 U7264 ( .AN(n5385), .B(n5384), .C(n5383), .Y(n5389) );
  AOI31X1 U7265 ( .A0(n5389), .A1(n5388), .A2(n5387), .B0(n5386), .Y(n5393) );
  AOI211X1 U7266 ( .A0(n5393), .A1(n5392), .B0(n5391), .C0(n5390), .Y(n5395)
         );
  AO21X1 U7267 ( .A0(cmd_valid), .A1(\state_cs[0] ), .B0(IRAM_valid), .Y(
        state_ns[1]) );
  NAND2X1 U7268 ( .A(n5399), .B(n5400), .Y(state_ns[0]) );
  NAND2X1 U7269 ( .A(cmd_valid), .B(n5403), .Y(n5402) );
  NAND4BX1 U7270 ( .AN(cmd[3]), .B(n5404), .C(n5405), .D(n5406), .Y(n5403) );
  OAI222XL U7271 ( .A0(n5415), .A1(n4953), .B0(n5416), .B1(n4956), .C0(n5418), 
        .C1(n5419), .Y(n5413) );
  OAI222XL U7272 ( .A0(n5426), .A1(n4952), .B0(n5427), .B1(n4956), .C0(n5428), 
        .C1(n4959), .Y(n5425) );
  MXI2X1 U7273 ( .A(\ImageBuffer[61][7] ), .B(n4949), .S0(n4875), .Y(n5431) );
  OAI222XL U7274 ( .A0(n5435), .A1(n4951), .B0(n5436), .B1(n4956), .C0(n5437), 
        .C1(n4958), .Y(n5434) );
  OAI222XL U7275 ( .A0(n5444), .A1(n4951), .B0(n5445), .B1(n4956), .C0(n5446), 
        .C1(n5419), .Y(n5443) );
  OAI222XL U7276 ( .A0(n5453), .A1(n4953), .B0(n5454), .B1(n4955), .C0(n5455), 
        .C1(n4959), .Y(n5452) );
  OAI222XL U7277 ( .A0(n5462), .A1(n4953), .B0(n5463), .B1(n4956), .C0(n5464), 
        .C1(n4959), .Y(n5461) );
  OAI222XL U7278 ( .A0(n5471), .A1(n4953), .B0(n5472), .B1(n4954), .C0(n5473), 
        .C1(n4959), .Y(n5470) );
  OAI222XL U7279 ( .A0(n5480), .A1(n4953), .B0(n5481), .B1(n4954), .C0(n5482), 
        .C1(n4959), .Y(n5479) );
  OAI222XL U7280 ( .A0(n5489), .A1(n4953), .B0(n5490), .B1(n5417), .C0(n5491), 
        .C1(n4959), .Y(n5488) );
  OAI222XL U7281 ( .A0(n5498), .A1(n4953), .B0(n5499), .B1(n4954), .C0(n5500), 
        .C1(n4959), .Y(n5497) );
  OAI222XL U7282 ( .A0(n5507), .A1(n4953), .B0(n5508), .B1(n5417), .C0(n5509), 
        .C1(n4959), .Y(n5506) );
  OAI222XL U7283 ( .A0(n5516), .A1(n4953), .B0(n5517), .B1(n4956), .C0(n5518), 
        .C1(n4959), .Y(n5515) );
  OAI222XL U7284 ( .A0(n5525), .A1(n4953), .B0(n5526), .B1(n4955), .C0(n5527), 
        .C1(n4959), .Y(n5524) );
  OAI222XL U7285 ( .A0(n5534), .A1(n4953), .B0(n5535), .B1(n5417), .C0(n5536), 
        .C1(n4959), .Y(n5533) );
  OAI222XL U7286 ( .A0(n5543), .A1(n4953), .B0(n5544), .B1(n5417), .C0(n5545), 
        .C1(n4959), .Y(n5542) );
  OAI222XL U7287 ( .A0(n5552), .A1(n4953), .B0(n5553), .B1(n4956), .C0(n5554), 
        .C1(n4959), .Y(n5551) );
  OAI222XL U7288 ( .A0(n5561), .A1(n4952), .B0(n5562), .B1(n4956), .C0(n5563), 
        .C1(n4958), .Y(n5560) );
  MXI2X1 U7289 ( .A(\ImageBuffer[46][7] ), .B(n4950), .S0(n4892), .Y(n5566) );
  AOI211X1 U7290 ( .A0(n5100), .A1(n5568), .B0(n5569), .C0(n5414), .Y(n5564)
         );
  OAI222XL U7291 ( .A0(n5570), .A1(n4952), .B0(n5571), .B1(n4956), .C0(n5572), 
        .C1(n4958), .Y(n5569) );
  OAI222XL U7292 ( .A0(n5579), .A1(n4952), .B0(n5580), .B1(n4956), .C0(n5581), 
        .C1(n4958), .Y(n5578) );
  MXI2X1 U7293 ( .A(\ImageBuffer[44][7] ), .B(n4950), .S0(n4894), .Y(n5584) );
  OAI222XL U7294 ( .A0(n5588), .A1(n4952), .B0(n5589), .B1(n4956), .C0(n5590), 
        .C1(n4958), .Y(n5587) );
  MXI2X1 U7295 ( .A(\ImageBuffer[43][7] ), .B(n4950), .S0(n4895), .Y(n5593) );
  OAI222XL U7296 ( .A0(n5597), .A1(n4952), .B0(n5598), .B1(n4956), .C0(n5599), 
        .C1(n4958), .Y(n5596) );
  OAI222XL U7297 ( .A0(n5606), .A1(n4952), .B0(n5607), .B1(n4956), .C0(n5608), 
        .C1(n4958), .Y(n5605) );
  MXI2X1 U7298 ( .A(\ImageBuffer[41][7] ), .B(n4950), .S0(n4897), .Y(n5611) );
  OAI222XL U7299 ( .A0(n5615), .A1(n4952), .B0(n5616), .B1(n4956), .C0(n5617), 
        .C1(n4958), .Y(n5614) );
  OAI222XL U7300 ( .A0(n5624), .A1(n4952), .B0(n5625), .B1(n4956), .C0(n5626), 
        .C1(n4958), .Y(n5623) );
  OAI222XL U7301 ( .A0(n5633), .A1(n4952), .B0(n5634), .B1(n4956), .C0(n5635), 
        .C1(n4958), .Y(n5632) );
  OAI222XL U7302 ( .A0(n5642), .A1(n4952), .B0(n5643), .B1(n4956), .C0(n5644), 
        .C1(n4958), .Y(n5641) );
  OAI222XL U7303 ( .A0(n5651), .A1(n4952), .B0(n5652), .B1(n4956), .C0(n5653), 
        .C1(n4958), .Y(n5650) );
  MXI2X1 U7304 ( .A(\ImageBuffer[36][7] ), .B(n4950), .S0(n4903), .Y(n5656) );
  OAI222XL U7305 ( .A0(n5660), .A1(n4952), .B0(n5661), .B1(n4956), .C0(n5662), 
        .C1(n4958), .Y(n5659) );
  OAI222XL U7306 ( .A0(n5669), .A1(n4951), .B0(n5670), .B1(n4955), .C0(n5671), 
        .C1(n5419), .Y(n5668) );
  OAI222XL U7307 ( .A0(n5678), .A1(n4951), .B0(n5679), .B1(n4955), .C0(n5680), 
        .C1(n4958), .Y(n5677) );
  OAI222XL U7308 ( .A0(n5687), .A1(n4951), .B0(n5688), .B1(n4955), .C0(n5689), 
        .C1(n5157), .Y(n5686) );
  OAI222XL U7309 ( .A0(n5696), .A1(n4951), .B0(n5697), .B1(n4955), .C0(n5698), 
        .C1(n4959), .Y(n5695) );
  OAI222XL U7310 ( .A0(n5705), .A1(n4951), .B0(n5706), .B1(n4955), .C0(n5707), 
        .C1(n4958), .Y(n5704) );
  OAI222XL U7311 ( .A0(n5714), .A1(n4951), .B0(n5715), .B1(n4955), .C0(n5716), 
        .C1(n5419), .Y(n5713) );
  OAI222XL U7312 ( .A0(n5723), .A1(n4951), .B0(n5724), .B1(n4955), .C0(n5725), 
        .C1(n4957), .Y(n5722) );
  OAI222XL U7313 ( .A0(n5732), .A1(n4951), .B0(n5733), .B1(n4955), .C0(n5734), 
        .C1(n4958), .Y(n5731) );
  OAI222XL U7314 ( .A0(n5741), .A1(n4951), .B0(n5742), .B1(n4955), .C0(n5743), 
        .C1(n5188), .Y(n5740) );
  OAI222XL U7315 ( .A0(n5750), .A1(n4951), .B0(n5751), .B1(n4955), .C0(n5752), 
        .C1(n4958), .Y(n5749) );
  OAI222XL U7316 ( .A0(n5759), .A1(n4951), .B0(n5760), .B1(n4955), .C0(n5761), 
        .C1(n4957), .Y(n5758) );
  OAI222XL U7317 ( .A0(n5768), .A1(n4951), .B0(n5769), .B1(n4955), .C0(n5770), 
        .C1(n4957), .Y(n5767) );
  OAI222XL U7318 ( .A0(n5777), .A1(n4951), .B0(n5778), .B1(n4954), .C0(n5779), 
        .C1(n4959), .Y(n5776) );
  OAI222XL U7319 ( .A0(n5786), .A1(n4951), .B0(n5787), .B1(n4954), .C0(n5788), 
        .C1(n4959), .Y(n5785) );
  OAI222XL U7320 ( .A0(n5795), .A1(n4951), .B0(n5796), .B1(n4954), .C0(n5797), 
        .C1(n4959), .Y(n5794) );
  OAI222XL U7321 ( .A0(n5804), .A1(n4952), .B0(n5805), .B1(n4954), .C0(n5806), 
        .C1(n4958), .Y(n5803) );
  OAI222XL U7322 ( .A0(n5813), .A1(n5310), .B0(n5814), .B1(n4954), .C0(n5815), 
        .C1(n4958), .Y(n5812) );
  OAI222XL U7323 ( .A0(n5822), .A1(n4951), .B0(n5823), .B1(n4954), .C0(n5824), 
        .C1(n4959), .Y(n5821) );
  OAI222XL U7324 ( .A0(n5831), .A1(n4951), .B0(n5832), .B1(n4954), .C0(n5833), 
        .C1(n4959), .Y(n5830) );
  MXI2X1 U7325 ( .A(\ImageBuffer[16][7] ), .B(n4948), .S0(n4925), .Y(n5836) );
  OAI222XL U7326 ( .A0(n5840), .A1(n5310), .B0(n5841), .B1(n4954), .C0(n5842), 
        .C1(n4957), .Y(n5839) );
  OAI222XL U7327 ( .A0(n5849), .A1(n4951), .B0(n5850), .B1(n4954), .C0(n5851), 
        .C1(n4959), .Y(n5848) );
  OAI222XL U7328 ( .A0(n5858), .A1(n4953), .B0(n5859), .B1(n4954), .C0(n5860), 
        .C1(n4957), .Y(n5857) );
  OAI222XL U7329 ( .A0(n5867), .A1(n4951), .B0(n5868), .B1(n4954), .C0(n5869), 
        .C1(n4959), .Y(n5866) );
  OAI222XL U7330 ( .A0(n5876), .A1(n5310), .B0(n5877), .B1(n4954), .C0(n5878), 
        .C1(n4957), .Y(n5875) );
  MXI2X1 U7331 ( .A(\ImageBuffer[11][7] ), .B(n4948), .S0(n4931), .Y(n5881) );
  OAI222XL U7332 ( .A0(n5885), .A1(n4952), .B0(n5886), .B1(n4955), .C0(n5887), 
        .C1(n4957), .Y(n5884) );
  MXI2X1 U7333 ( .A(\ImageBuffer[10][7] ), .B(n5410), .S0(n4932), .Y(n5890) );
  OAI222XL U7334 ( .A0(n5894), .A1(n4952), .B0(n5895), .B1(n4954), .C0(n5896), 
        .C1(n4957), .Y(n5893) );
  MXI2X1 U7335 ( .A(\ImageBuffer[9][7] ), .B(n5410), .S0(n4933), .Y(n5899) );
  OAI222XL U7336 ( .A0(n5903), .A1(n4952), .B0(n5904), .B1(n4954), .C0(n5905), 
        .C1(n4957), .Y(n5902) );
  MXI2X1 U7337 ( .A(\ImageBuffer[8][7] ), .B(n4949), .S0(n4934), .Y(n5908) );
  OAI222XL U7338 ( .A0(n5912), .A1(n4952), .B0(n5913), .B1(n4954), .C0(n5914), 
        .C1(n4957), .Y(n5911) );
  MXI2X1 U7339 ( .A(\ImageBuffer[7][7] ), .B(n4950), .S0(n4935), .Y(n5917) );
  OAI222XL U7340 ( .A0(n5921), .A1(n4953), .B0(n5922), .B1(n4955), .C0(n5923), 
        .C1(n4957), .Y(n5920) );
  MXI2X1 U7341 ( .A(\ImageBuffer[6][7] ), .B(n4948), .S0(n4936), .Y(n5926) );
  OAI222XL U7342 ( .A0(n5930), .A1(n4953), .B0(n5931), .B1(n4954), .C0(n5932), 
        .C1(n4957), .Y(n5929) );
  MXI2X1 U7343 ( .A(\ImageBuffer[5][7] ), .B(n4949), .S0(n4937), .Y(n5935) );
  OAI222XL U7344 ( .A0(n5939), .A1(n4953), .B0(n5940), .B1(n4955), .C0(n5941), 
        .C1(n4957), .Y(n5938) );
  MXI2X1 U7345 ( .A(\ImageBuffer[4][7] ), .B(n4950), .S0(n4938), .Y(n5944) );
  OAI222XL U7346 ( .A0(n5948), .A1(n4953), .B0(n5949), .B1(n4955), .C0(n5950), 
        .C1(n4957), .Y(n5947) );
  MXI2X1 U7347 ( .A(\ImageBuffer[3][7] ), .B(n4948), .S0(n4939), .Y(n5953) );
  OAI222XL U7348 ( .A0(n5957), .A1(n4953), .B0(n5958), .B1(n4954), .C0(n5959), 
        .C1(n4957), .Y(n5956) );
  MXI2X1 U7349 ( .A(\ImageBuffer[2][7] ), .B(n4949), .S0(n4940), .Y(n5962) );
  OAI222XL U7350 ( .A0(n5966), .A1(n4953), .B0(n5967), .B1(n4955), .C0(n5968), 
        .C1(n4957), .Y(n5965) );
  MXI2X1 U7351 ( .A(\ImageBuffer[1][7] ), .B(n4950), .S0(n4941), .Y(n5971) );
  OAI222XL U7352 ( .A0(n5975), .A1(n4953), .B0(n5976), .B1(n4956), .C0(n5977), 
        .C1(n4957), .Y(n5974) );
  MXI2X1 U7353 ( .A(\ImageBuffer[0][7] ), .B(n4950), .S0(n4942), .Y(n5980) );
  NOR2BX1 U7354 ( .AN(IROM_Q[7]), .B(n4945), .Y(n5410) );
  OAI222XL U7355 ( .A0(n5989), .A1(n4952), .B0(n5990), .B1(n4955), .C0(n5991), 
        .C1(n4957), .Y(n5984) );
  CLKINVX1 U7356 ( .A(n4861), .Y(n5419) );
  CLKINVX1 U7357 ( .A(N2766), .Y(n5417) );
  OAI222XL U7358 ( .A0(n5415), .A1(n4966), .B0(n5416), .B1(n4967), .C0(n5418), 
        .C1(n4973), .Y(n5995) );
  OAI222XL U7359 ( .A0(n5426), .A1(n4964), .B0(n5427), .B1(n5997), .C0(n5428), 
        .C1(n4971), .Y(n6000) );
  MXI2X1 U7360 ( .A(\ImageBuffer[61][6] ), .B(n4960), .S0(n4875), .Y(n6002) );
  OAI222XL U7361 ( .A0(n5435), .A1(n4966), .B0(n5436), .B1(n4969), .C0(n5437), 
        .C1(n4972), .Y(n6003) );
  OAI222XL U7362 ( .A0(n5444), .A1(n4963), .B0(n5445), .B1(n4968), .C0(n5446), 
        .C1(n4970), .Y(n6006) );
  OAI222XL U7363 ( .A0(n5453), .A1(n4966), .B0(n5454), .B1(n4969), .C0(n5455), 
        .C1(n4973), .Y(n6009) );
  MXI2X1 U7364 ( .A(\ImageBuffer[58][6] ), .B(n4962), .S0(n4878), .Y(n6011) );
  OAI222XL U7365 ( .A0(n5462), .A1(n4966), .B0(n5463), .B1(n4969), .C0(n5464), 
        .C1(n4973), .Y(n6012) );
  OAI222XL U7366 ( .A0(n5471), .A1(n4966), .B0(n5472), .B1(n4969), .C0(n5473), 
        .C1(n4973), .Y(n6015) );
  MXI2X1 U7367 ( .A(\ImageBuffer[56][6] ), .B(n4962), .S0(n4880), .Y(n6017) );
  OAI222XL U7368 ( .A0(n5480), .A1(n4966), .B0(n5481), .B1(n4969), .C0(n5482), 
        .C1(n4973), .Y(n6018) );
  OAI222XL U7369 ( .A0(n5489), .A1(n4966), .B0(n5490), .B1(n4969), .C0(n5491), 
        .C1(n4973), .Y(n6021) );
  MXI2X1 U7370 ( .A(\ImageBuffer[53][6] ), .B(n4962), .S0(n4884), .Y(n6026) );
  OAI222XL U7371 ( .A0(n5507), .A1(n4966), .B0(n5508), .B1(n4969), .C0(n5509), 
        .C1(n4973), .Y(n6027) );
  OAI222XL U7372 ( .A0(n5516), .A1(n4966), .B0(n5517), .B1(n4969), .C0(n5518), 
        .C1(n4973), .Y(n6030) );
  OAI222XL U7373 ( .A0(n5525), .A1(n4964), .B0(n5526), .B1(n4969), .C0(n5527), 
        .C1(n4973), .Y(n6033) );
  MXI2X1 U7374 ( .A(\ImageBuffer[50][6] ), .B(n4962), .S0(n4887), .Y(n6035) );
  OAI222XL U7375 ( .A0(n5534), .A1(n4966), .B0(n5535), .B1(n4969), .C0(n5536), 
        .C1(n4973), .Y(n6036) );
  OAI222XL U7376 ( .A0(n5543), .A1(n4966), .B0(n5544), .B1(n4969), .C0(n5545), 
        .C1(n4973), .Y(n6039) );
  OAI222XL U7377 ( .A0(n5552), .A1(n4965), .B0(n5553), .B1(n4969), .C0(n5554), 
        .C1(n4973), .Y(n6042) );
  OAI222XL U7378 ( .A0(n5561), .A1(n4965), .B0(n5562), .B1(n4967), .C0(n5563), 
        .C1(n4971), .Y(n6045) );
  MXI2X1 U7379 ( .A(\ImageBuffer[46][6] ), .B(n4961), .S0(n4892), .Y(n6047) );
  OAI222XL U7380 ( .A0(n5570), .A1(n4965), .B0(n5571), .B1(n5997), .C0(n5572), 
        .C1(n4971), .Y(n6048) );
  OAI222XL U7381 ( .A0(n5579), .A1(n4965), .B0(n5580), .B1(n4968), .C0(n5581), 
        .C1(n4973), .Y(n6051) );
  MXI2X1 U7382 ( .A(\ImageBuffer[44][6] ), .B(n4961), .S0(n4894), .Y(n6053) );
  OAI222XL U7383 ( .A0(n5588), .A1(n4965), .B0(n5589), .B1(n4968), .C0(n5590), 
        .C1(n4971), .Y(n6054) );
  OAI222XL U7384 ( .A0(n5597), .A1(n4965), .B0(n5598), .B1(n4967), .C0(n5599), 
        .C1(n4972), .Y(n6057) );
  OAI222XL U7385 ( .A0(n5606), .A1(n4965), .B0(n5607), .B1(n4969), .C0(n5608), 
        .C1(n4970), .Y(n6060) );
  MXI2X1 U7386 ( .A(\ImageBuffer[41][6] ), .B(n4961), .S0(n4897), .Y(n6062) );
  OAI222XL U7387 ( .A0(n5615), .A1(n4965), .B0(n5616), .B1(n4969), .C0(n5617), 
        .C1(n4971), .Y(n6063) );
  OAI222XL U7388 ( .A0(n5624), .A1(n4965), .B0(n5625), .B1(n4968), .C0(n5626), 
        .C1(n4973), .Y(n6066) );
  OAI222XL U7389 ( .A0(n5633), .A1(n4965), .B0(n5634), .B1(n4967), .C0(n5635), 
        .C1(n4970), .Y(n6069) );
  OAI222XL U7390 ( .A0(n5642), .A1(n4965), .B0(n5643), .B1(n4967), .C0(n5644), 
        .C1(n4972), .Y(n6072) );
  OAI222XL U7391 ( .A0(n5651), .A1(n4965), .B0(n5652), .B1(n4969), .C0(n5653), 
        .C1(n4973), .Y(n6075) );
  MXI2X1 U7392 ( .A(\ImageBuffer[36][6] ), .B(n4961), .S0(n4903), .Y(n6077) );
  OAI222XL U7393 ( .A0(n5660), .A1(n4965), .B0(n5661), .B1(n4968), .C0(n5662), 
        .C1(n4971), .Y(n6078) );
  OAI222XL U7394 ( .A0(n5669), .A1(n4966), .B0(n5670), .B1(n4968), .C0(n5671), 
        .C1(n4972), .Y(n6081) );
  OAI222XL U7395 ( .A0(n5678), .A1(n4966), .B0(n5679), .B1(n4969), .C0(n5680), 
        .C1(n4972), .Y(n6084) );
  OAI222XL U7396 ( .A0(n5687), .A1(n4966), .B0(n5688), .B1(n4967), .C0(n5689), 
        .C1(n4972), .Y(n6087) );
  OAI222XL U7397 ( .A0(n5696), .A1(n4965), .B0(n5697), .B1(n4968), .C0(n5698), 
        .C1(n4972), .Y(n6090) );
  OAI222XL U7398 ( .A0(n5705), .A1(n4964), .B0(n5706), .B1(n4967), .C0(n5707), 
        .C1(n4972), .Y(n6093) );
  OAI222XL U7399 ( .A0(n5714), .A1(n4963), .B0(n5715), .B1(n4969), .C0(n5716), 
        .C1(n4972), .Y(n6096) );
  OAI222XL U7400 ( .A0(n5723), .A1(n4963), .B0(n5724), .B1(n4969), .C0(n5725), 
        .C1(n4972), .Y(n6099) );
  OAI222XL U7401 ( .A0(n5732), .A1(n4965), .B0(n5733), .B1(n4968), .C0(n5734), 
        .C1(n4972), .Y(n6102) );
  OAI222XL U7402 ( .A0(n5741), .A1(n4966), .B0(n5742), .B1(n4967), .C0(n5743), 
        .C1(n4972), .Y(n6105) );
  OAI222XL U7403 ( .A0(n5750), .A1(n4966), .B0(n5751), .B1(n5997), .C0(n5752), 
        .C1(n4972), .Y(n6108) );
  OAI222XL U7404 ( .A0(n5759), .A1(n4966), .B0(n5760), .B1(n4969), .C0(n5761), 
        .C1(n4972), .Y(n6111) );
  OAI222XL U7405 ( .A0(n5768), .A1(n4966), .B0(n5769), .B1(n5997), .C0(n5770), 
        .C1(n4972), .Y(n6114) );
  OAI222XL U7406 ( .A0(n5777), .A1(n4964), .B0(n5778), .B1(n4968), .C0(n5779), 
        .C1(n4971), .Y(n6117) );
  OAI222XL U7407 ( .A0(n5786), .A1(n4964), .B0(n5787), .B1(n4968), .C0(n5788), 
        .C1(n4971), .Y(n6120) );
  OAI222XL U7408 ( .A0(n5795), .A1(n4964), .B0(n5796), .B1(n4968), .C0(n5797), 
        .C1(n4971), .Y(n6123) );
  OAI222XL U7409 ( .A0(n5804), .A1(n4964), .B0(n5805), .B1(n4968), .C0(n5806), 
        .C1(n4971), .Y(n6126) );
  MXI2X1 U7410 ( .A(\ImageBuffer[19][6] ), .B(n4960), .S0(n4922), .Y(n6128) );
  OAI222XL U7411 ( .A0(n5813), .A1(n4964), .B0(n5814), .B1(n4968), .C0(n5815), 
        .C1(n4971), .Y(n6129) );
  OAI222XL U7412 ( .A0(n5822), .A1(n4964), .B0(n5823), .B1(n4968), .C0(n5824), 
        .C1(n4971), .Y(n6132) );
  OAI222XL U7413 ( .A0(n5831), .A1(n4964), .B0(n5832), .B1(n4968), .C0(n5833), 
        .C1(n4971), .Y(n6135) );
  MXI2X1 U7414 ( .A(\ImageBuffer[16][6] ), .B(n4962), .S0(n4925), .Y(n6137) );
  OAI222XL U7415 ( .A0(n5840), .A1(n4964), .B0(n5841), .B1(n4968), .C0(n5842), 
        .C1(n4971), .Y(n6138) );
  OAI222XL U7416 ( .A0(n5849), .A1(n4964), .B0(n5850), .B1(n4968), .C0(n5851), 
        .C1(n4971), .Y(n6141) );
  OAI222XL U7417 ( .A0(n5858), .A1(n4964), .B0(n5859), .B1(n4968), .C0(n5860), 
        .C1(n4971), .Y(n6144) );
  OAI222XL U7418 ( .A0(n5867), .A1(n4964), .B0(n5868), .B1(n4968), .C0(n5869), 
        .C1(n4971), .Y(n6147) );
  OAI222XL U7419 ( .A0(n5876), .A1(n4964), .B0(n5877), .B1(n4968), .C0(n5878), 
        .C1(n4971), .Y(n6150) );
  MXI2X1 U7420 ( .A(\ImageBuffer[11][6] ), .B(n4962), .S0(n4931), .Y(n6152) );
  OAI222XL U7421 ( .A0(n5885), .A1(n4963), .B0(n5886), .B1(n4967), .C0(n5887), 
        .C1(n4970), .Y(n6153) );
  MXI2X1 U7422 ( .A(\ImageBuffer[10][6] ), .B(n4961), .S0(n4932), .Y(n6155) );
  OAI222XL U7423 ( .A0(n5894), .A1(n4963), .B0(n5895), .B1(n4967), .C0(n5896), 
        .C1(n4970), .Y(n6156) );
  MXI2X1 U7424 ( .A(\ImageBuffer[9][6] ), .B(n4960), .S0(n4933), .Y(n6158) );
  OAI222XL U7425 ( .A0(n5903), .A1(n4963), .B0(n5904), .B1(n4967), .C0(n5905), 
        .C1(n4970), .Y(n6159) );
  MXI2X1 U7426 ( .A(\ImageBuffer[8][6] ), .B(n4962), .S0(n4934), .Y(n6161) );
  OAI222XL U7427 ( .A0(n5912), .A1(n4963), .B0(n5913), .B1(n4967), .C0(n5914), 
        .C1(n4970), .Y(n6162) );
  MXI2X1 U7428 ( .A(\ImageBuffer[7][6] ), .B(n4961), .S0(n4935), .Y(n6164) );
  OAI222XL U7429 ( .A0(n5921), .A1(n4963), .B0(n5922), .B1(n4967), .C0(n5923), 
        .C1(n4970), .Y(n6165) );
  MXI2X1 U7430 ( .A(\ImageBuffer[6][6] ), .B(n4960), .S0(n4936), .Y(n6167) );
  OAI222XL U7431 ( .A0(n5930), .A1(n4963), .B0(n5931), .B1(n4967), .C0(n5932), 
        .C1(n4970), .Y(n6168) );
  MXI2X1 U7432 ( .A(\ImageBuffer[5][6] ), .B(n4962), .S0(n4937), .Y(n6170) );
  OAI222XL U7433 ( .A0(n5939), .A1(n4963), .B0(n5940), .B1(n4967), .C0(n5941), 
        .C1(n4970), .Y(n6171) );
  MXI2X1 U7434 ( .A(\ImageBuffer[4][6] ), .B(n4961), .S0(n4938), .Y(n6173) );
  OAI222XL U7435 ( .A0(n5948), .A1(n4963), .B0(n5949), .B1(n4967), .C0(n5950), 
        .C1(n4970), .Y(n6174) );
  MXI2X1 U7436 ( .A(\ImageBuffer[3][6] ), .B(n4960), .S0(n4939), .Y(n6176) );
  OAI222XL U7437 ( .A0(n5957), .A1(n4963), .B0(n5958), .B1(n4967), .C0(n5959), 
        .C1(n4970), .Y(n6177) );
  MXI2X1 U7438 ( .A(\ImageBuffer[2][6] ), .B(n5994), .S0(n4940), .Y(n6179) );
  MXI2X1 U7439 ( .A(\ImageBuffer[1][6] ), .B(n5994), .S0(n4941), .Y(n6182) );
  OAI222XL U7440 ( .A0(n5975), .A1(n4963), .B0(n5976), .B1(n4967), .C0(n5977), 
        .C1(n4970), .Y(n6183) );
  MXI2X1 U7441 ( .A(\ImageBuffer[0][6] ), .B(n4960), .S0(n4942), .Y(n6185) );
  NOR2BX1 U7442 ( .AN(IROM_Q[6]), .B(n4945), .Y(n5994) );
  OAI222XL U7443 ( .A0(n5989), .A1(n4963), .B0(n5990), .B1(n4967), .C0(n5991), 
        .C1(n4970), .Y(n6186) );
  CLKINVX1 U7444 ( .A(N2767), .Y(n5997) );
  OAI21XL U7445 ( .A0(n6188), .A1(n5408), .B0(n6189), .Y(n8218) );
  AOI211X1 U7446 ( .A0(n5092), .A1(n5412), .B0(n6191), .C0(n3349), .Y(n6188)
         );
  OAI222XL U7447 ( .A0(n5415), .A1(n4977), .B0(n5416), .B1(n4982), .C0(n5418), 
        .C1(n4984), .Y(n6191) );
  OAI21XL U7448 ( .A0(n6196), .A1(n5421), .B0(n6197), .Y(n8219) );
  AOI211X1 U7449 ( .A0(n5092), .A1(n5424), .B0(n6198), .C0(n6192), .Y(n6196)
         );
  OAI222XL U7450 ( .A0(n5426), .A1(n4979), .B0(n5427), .B1(n4982), .C0(n5428), 
        .C1(n4985), .Y(n6198) );
  OAI21XL U7451 ( .A0(n6199), .A1(n5430), .B0(n6200), .Y(n8220) );
  AOI211X1 U7452 ( .A0(n5092), .A1(n5433), .B0(n6201), .C0(n3350), .Y(n6199)
         );
  OAI21XL U7453 ( .A0(n6202), .A1(n5439), .B0(n6203), .Y(n8221) );
  AOI211X1 U7454 ( .A0(n5092), .A1(n5442), .B0(n6204), .C0(n6192), .Y(n6202)
         );
  OAI222XL U7455 ( .A0(n5444), .A1(n4979), .B0(n5445), .B1(n4982), .C0(n5446), 
        .C1(n4984), .Y(n6204) );
  OAI21XL U7456 ( .A0(n6205), .A1(n5448), .B0(n6206), .Y(n8222) );
  AOI211X1 U7457 ( .A0(n5092), .A1(n5451), .B0(n6207), .C0(n3350), .Y(n6205)
         );
  OAI222XL U7458 ( .A0(n5453), .A1(n4979), .B0(n5454), .B1(n4982), .C0(n5455), 
        .C1(n4985), .Y(n6207) );
  OAI21XL U7459 ( .A0(n6208), .A1(n5457), .B0(n6209), .Y(n8223) );
  MXI2X1 U7460 ( .A(\ImageBuffer[58][5] ), .B(n4976), .S0(n4878), .Y(n6209) );
  AOI211X1 U7461 ( .A0(n5092), .A1(n5460), .B0(n6210), .C0(n3349), .Y(n6208)
         );
  OAI222XL U7462 ( .A0(n5462), .A1(n4979), .B0(n5463), .B1(n4981), .C0(n5464), 
        .C1(n4985), .Y(n6210) );
  OAI21XL U7463 ( .A0(n6211), .A1(n5466), .B0(n6212), .Y(n8224) );
  AOI211X1 U7464 ( .A0(n5092), .A1(n5469), .B0(n6213), .C0(n6192), .Y(n6211)
         );
  OAI222XL U7465 ( .A0(n5471), .A1(n4979), .B0(n5472), .B1(n4982), .C0(n5473), 
        .C1(n6195), .Y(n6213) );
  OAI21XL U7466 ( .A0(n6214), .A1(n5475), .B0(n6215), .Y(n8225) );
  MXI2X1 U7467 ( .A(\ImageBuffer[56][5] ), .B(n4976), .S0(n4880), .Y(n6215) );
  AOI211X1 U7468 ( .A0(n5092), .A1(n5478), .B0(n6216), .C0(n3350), .Y(n6214)
         );
  OAI222XL U7469 ( .A0(n5480), .A1(n4979), .B0(n5481), .B1(n4982), .C0(n5482), 
        .C1(n4983), .Y(n6216) );
  OAI21XL U7470 ( .A0(n6217), .A1(n5484), .B0(n6218), .Y(n8226) );
  AOI211X1 U7471 ( .A0(n5092), .A1(n5487), .B0(n6219), .C0(n3349), .Y(n6217)
         );
  OAI222XL U7472 ( .A0(n5489), .A1(n4979), .B0(n5490), .B1(n4982), .C0(n5491), 
        .C1(n4983), .Y(n6219) );
  OAI21XL U7473 ( .A0(n6220), .A1(n5493), .B0(n6221), .Y(n8227) );
  AOI211X1 U7474 ( .A0(n5092), .A1(n5496), .B0(n6222), .C0(n3350), .Y(n6220)
         );
  OAI21XL U7475 ( .A0(n6223), .A1(n5502), .B0(n6224), .Y(n8228) );
  AOI211X1 U7476 ( .A0(n5092), .A1(n5505), .B0(n6225), .C0(n6192), .Y(n6223)
         );
  OAI222XL U7477 ( .A0(n5507), .A1(n4979), .B0(n5508), .B1(n4982), .C0(n5509), 
        .C1(n6195), .Y(n6225) );
  OAI21XL U7478 ( .A0(n6226), .A1(n5511), .B0(n6227), .Y(n8229) );
  AOI211X1 U7479 ( .A0(n5092), .A1(n5514), .B0(n6228), .C0(n3349), .Y(n6226)
         );
  OAI222XL U7480 ( .A0(n5516), .A1(n4979), .B0(n5517), .B1(n4982), .C0(n5518), 
        .C1(n4984), .Y(n6228) );
  OAI21XL U7481 ( .A0(n6229), .A1(n5520), .B0(n6230), .Y(n8230) );
  AOI211X1 U7482 ( .A0(n5092), .A1(n5523), .B0(n6231), .C0(n3350), .Y(n6229)
         );
  OAI222XL U7483 ( .A0(n5525), .A1(n4979), .B0(n5526), .B1(n4982), .C0(n5527), 
        .C1(n4983), .Y(n6231) );
  OAI21XL U7484 ( .A0(n6232), .A1(n5529), .B0(n6233), .Y(n8231) );
  MXI2X1 U7485 ( .A(\ImageBuffer[50][5] ), .B(n4976), .S0(n4887), .Y(n6233) );
  AOI211X1 U7486 ( .A0(n5092), .A1(n5532), .B0(n6234), .C0(n3349), .Y(n6232)
         );
  OAI222XL U7487 ( .A0(n5534), .A1(n4979), .B0(n5535), .B1(n4982), .C0(n5536), 
        .C1(n6195), .Y(n6234) );
  OAI21XL U7488 ( .A0(n6235), .A1(n5538), .B0(n6236), .Y(n8232) );
  AOI211X1 U7489 ( .A0(n5092), .A1(n5541), .B0(n6237), .C0(n6192), .Y(n6235)
         );
  OAI222XL U7490 ( .A0(n5543), .A1(n4979), .B0(n5544), .B1(n4982), .C0(n5545), 
        .C1(n6195), .Y(n6237) );
  OAI21XL U7491 ( .A0(n6238), .A1(n5547), .B0(n6239), .Y(n8233) );
  AOI211X1 U7492 ( .A0(n5092), .A1(n5550), .B0(n6240), .C0(n3349), .Y(n6238)
         );
  OAI222XL U7493 ( .A0(n5552), .A1(n4979), .B0(n5553), .B1(n4981), .C0(n5554), 
        .C1(n4985), .Y(n6240) );
  OAI21XL U7494 ( .A0(n6241), .A1(n5556), .B0(n6242), .Y(n8234) );
  AOI211X1 U7495 ( .A0(n3361), .A1(n5559), .B0(n6243), .C0(n6192), .Y(n6241)
         );
  OAI222XL U7496 ( .A0(n5561), .A1(n4978), .B0(n5562), .B1(n4981), .C0(n5563), 
        .C1(n4985), .Y(n6243) );
  OAI21XL U7497 ( .A0(n6244), .A1(n5565), .B0(n6245), .Y(n8235) );
  MXI2X1 U7498 ( .A(\ImageBuffer[46][5] ), .B(n4975), .S0(n4892), .Y(n6245) );
  AOI211X1 U7499 ( .A0(n5092), .A1(n5568), .B0(n6246), .C0(n6192), .Y(n6244)
         );
  OAI222XL U7500 ( .A0(n5570), .A1(n4978), .B0(n5571), .B1(n4981), .C0(n5572), 
        .C1(n4984), .Y(n6246) );
  OAI21XL U7501 ( .A0(n6247), .A1(n5574), .B0(n6248), .Y(n8236) );
  AOI211X1 U7502 ( .A0(n5093), .A1(n5577), .B0(n6249), .C0(n3350), .Y(n6247)
         );
  OAI222XL U7503 ( .A0(n5579), .A1(n4978), .B0(n5580), .B1(n4981), .C0(n5581), 
        .C1(n4984), .Y(n6249) );
  OAI21XL U7504 ( .A0(n6250), .A1(n5583), .B0(n6251), .Y(n8237) );
  MXI2X1 U7505 ( .A(\ImageBuffer[44][5] ), .B(n4975), .S0(n4894), .Y(n6251) );
  AOI211X1 U7506 ( .A0(n5092), .A1(n5586), .B0(n6252), .C0(n3349), .Y(n6250)
         );
  OAI222XL U7507 ( .A0(n5588), .A1(n4978), .B0(n5589), .B1(n4981), .C0(n5590), 
        .C1(n4984), .Y(n6252) );
  OAI21XL U7508 ( .A0(n6253), .A1(n5592), .B0(n6254), .Y(n8238) );
  AOI211X1 U7509 ( .A0(n3361), .A1(n5595), .B0(n6255), .C0(n3349), .Y(n6253)
         );
  OAI222XL U7510 ( .A0(n5597), .A1(n4978), .B0(n5598), .B1(n4981), .C0(n5599), 
        .C1(n4985), .Y(n6255) );
  OAI21XL U7511 ( .A0(n6256), .A1(n5601), .B0(n6257), .Y(n8239) );
  AOI211X1 U7512 ( .A0(n5093), .A1(n5604), .B0(n6258), .C0(n6192), .Y(n6256)
         );
  OAI222XL U7513 ( .A0(n5606), .A1(n4978), .B0(n5607), .B1(n4981), .C0(n5608), 
        .C1(n4983), .Y(n6258) );
  OAI21XL U7514 ( .A0(n6259), .A1(n5610), .B0(n6260), .Y(n8240) );
  MXI2X1 U7515 ( .A(\ImageBuffer[41][5] ), .B(n4975), .S0(n4897), .Y(n6260) );
  AOI211X1 U7516 ( .A0(n5092), .A1(n5613), .B0(n6261), .C0(n6192), .Y(n6259)
         );
  OAI222XL U7517 ( .A0(n5615), .A1(n4978), .B0(n5616), .B1(n4981), .C0(n5617), 
        .C1(n4983), .Y(n6261) );
  OAI21XL U7518 ( .A0(n6262), .A1(n5619), .B0(n6263), .Y(n8241) );
  AOI211X1 U7519 ( .A0(n5092), .A1(n5622), .B0(n6264), .C0(n3350), .Y(n6262)
         );
  OAI222XL U7520 ( .A0(n5624), .A1(n4978), .B0(n5625), .B1(n4981), .C0(n5626), 
        .C1(n4985), .Y(n6264) );
  OAI21XL U7521 ( .A0(n6265), .A1(n5628), .B0(n6266), .Y(n8242) );
  AOI211X1 U7522 ( .A0(n3361), .A1(n5631), .B0(n6267), .C0(n3350), .Y(n6265)
         );
  OAI222XL U7523 ( .A0(n5633), .A1(n4978), .B0(n5634), .B1(n4981), .C0(n5635), 
        .C1(n4984), .Y(n6267) );
  OAI21XL U7524 ( .A0(n6268), .A1(n5637), .B0(n6269), .Y(n8243) );
  AOI211X1 U7525 ( .A0(n5093), .A1(n5640), .B0(n6270), .C0(n3349), .Y(n6268)
         );
  OAI222XL U7526 ( .A0(n5642), .A1(n4978), .B0(n5643), .B1(n4981), .C0(n5644), 
        .C1(n4984), .Y(n6270) );
  OAI21XL U7527 ( .A0(n6271), .A1(n5646), .B0(n6272), .Y(n8244) );
  AOI211X1 U7528 ( .A0(n3361), .A1(n5649), .B0(n6273), .C0(n6192), .Y(n6271)
         );
  OAI222XL U7529 ( .A0(n5651), .A1(n4978), .B0(n5652), .B1(n4981), .C0(n5653), 
        .C1(n4983), .Y(n6273) );
  OAI21XL U7530 ( .A0(n6274), .A1(n5655), .B0(n6275), .Y(n8245) );
  AOI211X1 U7531 ( .A0(n5093), .A1(n5658), .B0(n6276), .C0(n3350), .Y(n6274)
         );
  OAI222XL U7532 ( .A0(n5660), .A1(n4978), .B0(n5661), .B1(n4981), .C0(n5662), 
        .C1(n4985), .Y(n6276) );
  OAI21XL U7533 ( .A0(n6277), .A1(n5664), .B0(n6278), .Y(n8246) );
  AOI211X1 U7534 ( .A0(n5092), .A1(n5667), .B0(n6279), .C0(n3350), .Y(n6277)
         );
  OAI222XL U7535 ( .A0(n5669), .A1(n4977), .B0(n5670), .B1(n4980), .C0(n5671), 
        .C1(n4985), .Y(n6279) );
  OAI21XL U7536 ( .A0(n6280), .A1(n5673), .B0(n6281), .Y(n8247) );
  AOI211X1 U7537 ( .A0(n3361), .A1(n5676), .B0(n6282), .C0(n3350), .Y(n6280)
         );
  OAI222XL U7538 ( .A0(n5678), .A1(n4977), .B0(n5679), .B1(n4980), .C0(n5680), 
        .C1(n4985), .Y(n6282) );
  OAI21XL U7539 ( .A0(n6283), .A1(n5682), .B0(n6284), .Y(n8248) );
  AOI211X1 U7540 ( .A0(n5092), .A1(n5685), .B0(n6285), .C0(n6192), .Y(n6283)
         );
  OAI222XL U7541 ( .A0(n5687), .A1(n4977), .B0(n5688), .B1(n4981), .C0(n5689), 
        .C1(n4985), .Y(n6285) );
  OAI21XL U7542 ( .A0(n6286), .A1(n5691), .B0(n6287), .Y(n8249) );
  AOI211X1 U7543 ( .A0(n5092), .A1(n5694), .B0(n6288), .C0(n3349), .Y(n6286)
         );
  OAI222XL U7544 ( .A0(n5696), .A1(n4977), .B0(n5697), .B1(n6194), .C0(n5698), 
        .C1(n4985), .Y(n6288) );
  OAI21XL U7545 ( .A0(n6289), .A1(n5700), .B0(n6290), .Y(n8250) );
  AOI211X1 U7546 ( .A0(n5093), .A1(n5703), .B0(n6291), .C0(n3349), .Y(n6289)
         );
  OAI222XL U7547 ( .A0(n5705), .A1(n4977), .B0(n5706), .B1(n4981), .C0(n5707), 
        .C1(n4985), .Y(n6291) );
  OAI21XL U7548 ( .A0(n6292), .A1(n5709), .B0(n6293), .Y(n8251) );
  AOI211X1 U7549 ( .A0(n5092), .A1(n5712), .B0(n6294), .C0(n3350), .Y(n6292)
         );
  OAI222XL U7550 ( .A0(n5714), .A1(n4977), .B0(n5715), .B1(n4982), .C0(n5716), 
        .C1(n4985), .Y(n6294) );
  OAI21XL U7551 ( .A0(n6295), .A1(n5718), .B0(n6296), .Y(n8252) );
  AOI211X1 U7552 ( .A0(n5092), .A1(n5721), .B0(n6297), .C0(n6192), .Y(n6295)
         );
  OAI222XL U7553 ( .A0(n5723), .A1(n4977), .B0(n5724), .B1(n4982), .C0(n5725), 
        .C1(n4985), .Y(n6297) );
  OAI21XL U7554 ( .A0(n6298), .A1(n5727), .B0(n6299), .Y(n8253) );
  AOI211X1 U7555 ( .A0(n5092), .A1(n5730), .B0(n6300), .C0(n3349), .Y(n6298)
         );
  OAI222XL U7556 ( .A0(n5732), .A1(n4977), .B0(n5733), .B1(n4980), .C0(n5734), 
        .C1(n4985), .Y(n6300) );
  OAI21XL U7557 ( .A0(n6301), .A1(n5736), .B0(n6302), .Y(n8254) );
  AOI211X1 U7558 ( .A0(n3361), .A1(n5739), .B0(n6303), .C0(n6192), .Y(n6301)
         );
  OAI222XL U7559 ( .A0(n5741), .A1(n4977), .B0(n5742), .B1(n4980), .C0(n5743), 
        .C1(n4985), .Y(n6303) );
  OAI21XL U7560 ( .A0(n6304), .A1(n5745), .B0(n6305), .Y(n8255) );
  AOI211X1 U7561 ( .A0(n5093), .A1(n5748), .B0(n6306), .C0(n6192), .Y(n6304)
         );
  OAI222XL U7562 ( .A0(n5750), .A1(n4977), .B0(n5751), .B1(n4980), .C0(n5752), 
        .C1(n4985), .Y(n6306) );
  OAI21XL U7563 ( .A0(n6307), .A1(n5754), .B0(n6308), .Y(n8256) );
  AOI211X1 U7564 ( .A0(n3361), .A1(n5757), .B0(n6309), .C0(n3350), .Y(n6307)
         );
  OAI222XL U7565 ( .A0(n5759), .A1(n4977), .B0(n5760), .B1(n4981), .C0(n5761), 
        .C1(n4985), .Y(n6309) );
  OAI21XL U7566 ( .A0(n6310), .A1(n5763), .B0(n6311), .Y(n8257) );
  AOI211X1 U7567 ( .A0(n5093), .A1(n5766), .B0(n6312), .C0(n3349), .Y(n6310)
         );
  OAI222XL U7568 ( .A0(n5768), .A1(n4977), .B0(n5769), .B1(n4982), .C0(n5770), 
        .C1(n4985), .Y(n6312) );
  OAI21XL U7569 ( .A0(n6313), .A1(n5772), .B0(n6314), .Y(n8258) );
  AOI211X1 U7570 ( .A0(n3360), .A1(n5775), .B0(n6315), .C0(n3349), .Y(n6313)
         );
  OAI222XL U7571 ( .A0(n5777), .A1(n4977), .B0(n5778), .B1(n4980), .C0(n5779), 
        .C1(n4984), .Y(n6315) );
  OAI21XL U7572 ( .A0(n6316), .A1(n5781), .B0(n6317), .Y(n8259) );
  AOI211X1 U7573 ( .A0(n3361), .A1(n5784), .B0(n6318), .C0(n3350), .Y(n6316)
         );
  OAI222XL U7574 ( .A0(n5786), .A1(n4977), .B0(n5787), .B1(n4981), .C0(n5788), 
        .C1(n4984), .Y(n6318) );
  OAI21XL U7575 ( .A0(n6319), .A1(n5790), .B0(n6320), .Y(n8260) );
  AOI211X1 U7576 ( .A0(n5093), .A1(n5793), .B0(n6321), .C0(n6192), .Y(n6319)
         );
  OAI222XL U7577 ( .A0(n5795), .A1(n6193), .B0(n5796), .B1(n4982), .C0(n5797), 
        .C1(n4984), .Y(n6321) );
  OAI21XL U7578 ( .A0(n6322), .A1(n5799), .B0(n6323), .Y(n8261) );
  AOI211X1 U7579 ( .A0(n5092), .A1(n5802), .B0(n6324), .C0(n3349), .Y(n6322)
         );
  OAI222XL U7580 ( .A0(n5804), .A1(n4979), .B0(n5805), .B1(n4980), .C0(n5806), 
        .C1(n4984), .Y(n6324) );
  OAI21XL U7581 ( .A0(n6325), .A1(n5808), .B0(n6326), .Y(n8262) );
  MXI2X1 U7582 ( .A(\ImageBuffer[19][5] ), .B(n4974), .S0(n4922), .Y(n6326) );
  AOI211X1 U7583 ( .A0(n5092), .A1(n5811), .B0(n6327), .C0(n3349), .Y(n6325)
         );
  OAI222XL U7584 ( .A0(n5813), .A1(n4978), .B0(n5814), .B1(n4982), .C0(n5815), 
        .C1(n4984), .Y(n6327) );
  OAI21XL U7585 ( .A0(n6328), .A1(n5817), .B0(n6329), .Y(n8263) );
  AOI211X1 U7586 ( .A0(n3360), .A1(n5820), .B0(n6330), .C0(n3349), .Y(n6328)
         );
  OAI222XL U7587 ( .A0(n5822), .A1(n4978), .B0(n5823), .B1(n4982), .C0(n5824), 
        .C1(n4984), .Y(n6330) );
  OAI21XL U7588 ( .A0(n6331), .A1(n5826), .B0(n6332), .Y(n8264) );
  AOI211X1 U7589 ( .A0(n5092), .A1(n5829), .B0(n6333), .C0(n3350), .Y(n6331)
         );
  OAI21XL U7590 ( .A0(n6334), .A1(n5835), .B0(n6335), .Y(n8265) );
  MXI2X1 U7591 ( .A(\ImageBuffer[16][5] ), .B(n4976), .S0(n4925), .Y(n6335) );
  AOI211X1 U7592 ( .A0(n5092), .A1(n5838), .B0(n6336), .C0(n3350), .Y(n6334)
         );
  OAI222XL U7593 ( .A0(n5840), .A1(n4977), .B0(n5841), .B1(n4982), .C0(n5842), 
        .C1(n4984), .Y(n6336) );
  OAI21XL U7594 ( .A0(n6337), .A1(n5844), .B0(n6338), .Y(n8266) );
  AOI211X1 U7595 ( .A0(n5092), .A1(n5847), .B0(n6339), .C0(n6192), .Y(n6337)
         );
  OAI222XL U7596 ( .A0(n5849), .A1(n4979), .B0(n5850), .B1(n6194), .C0(n5851), 
        .C1(n4984), .Y(n6339) );
  OAI21XL U7597 ( .A0(n6340), .A1(n5853), .B0(n6341), .Y(n8267) );
  AOI211X1 U7598 ( .A0(n5093), .A1(n5856), .B0(n6342), .C0(n3350), .Y(n6340)
         );
  OAI222XL U7599 ( .A0(n5858), .A1(n4978), .B0(n5859), .B1(n6194), .C0(n5860), 
        .C1(n4984), .Y(n6342) );
  OAI21XL U7600 ( .A0(n6343), .A1(n5862), .B0(n6344), .Y(n8268) );
  AOI211X1 U7601 ( .A0(n5092), .A1(n5865), .B0(n6345), .C0(n3349), .Y(n6343)
         );
  OAI222XL U7602 ( .A0(n5867), .A1(n4977), .B0(n5868), .B1(n6194), .C0(n5869), 
        .C1(n4984), .Y(n6345) );
  OAI21XL U7603 ( .A0(n6346), .A1(n5871), .B0(n6347), .Y(n8269) );
  AOI211X1 U7604 ( .A0(n3361), .A1(n5874), .B0(n6348), .C0(n6192), .Y(n6346)
         );
  OAI222XL U7605 ( .A0(n5876), .A1(n4978), .B0(n5877), .B1(n4981), .C0(n5878), 
        .C1(n4984), .Y(n6348) );
  OAI21XL U7606 ( .A0(n6349), .A1(n5880), .B0(n6350), .Y(n8270) );
  MXI2X1 U7607 ( .A(\ImageBuffer[11][5] ), .B(n4975), .S0(n4931), .Y(n6350) );
  AOI211X1 U7608 ( .A0(n5092), .A1(n5883), .B0(n6351), .C0(n6192), .Y(n6349)
         );
  OAI222XL U7609 ( .A0(n5885), .A1(n4978), .B0(n5886), .B1(n4980), .C0(n5887), 
        .C1(n4983), .Y(n6351) );
  OAI21XL U7610 ( .A0(n6352), .A1(n5889), .B0(n6353), .Y(n8271) );
  MXI2X1 U7611 ( .A(\ImageBuffer[10][5] ), .B(n4974), .S0(n4932), .Y(n6353) );
  AOI211X1 U7612 ( .A0(n5092), .A1(n5892), .B0(n6354), .C0(n3350), .Y(n6352)
         );
  OAI222XL U7613 ( .A0(n5894), .A1(n4977), .B0(n5895), .B1(n4980), .C0(n5896), 
        .C1(n4983), .Y(n6354) );
  OAI21XL U7614 ( .A0(n6355), .A1(n5898), .B0(n6356), .Y(n8272) );
  MXI2X1 U7615 ( .A(\ImageBuffer[9][5] ), .B(n4976), .S0(n4933), .Y(n6356) );
  AOI211X1 U7616 ( .A0(n5092), .A1(n5901), .B0(n6357), .C0(n3349), .Y(n6355)
         );
  OAI222XL U7617 ( .A0(n5903), .A1(n4977), .B0(n5904), .B1(n4980), .C0(n5905), 
        .C1(n4983), .Y(n6357) );
  OAI21XL U7618 ( .A0(n6358), .A1(n5907), .B0(n6359), .Y(n8273) );
  MXI2X1 U7619 ( .A(\ImageBuffer[8][5] ), .B(n4975), .S0(n4934), .Y(n6359) );
  AOI211X1 U7620 ( .A0(n5092), .A1(n5910), .B0(n6360), .C0(n6192), .Y(n6358)
         );
  OAI222XL U7621 ( .A0(n5912), .A1(n6193), .B0(n5913), .B1(n4980), .C0(n5914), 
        .C1(n4983), .Y(n6360) );
  OAI21XL U7622 ( .A0(n6361), .A1(n5916), .B0(n6362), .Y(n8274) );
  MXI2X1 U7623 ( .A(\ImageBuffer[7][5] ), .B(n4974), .S0(n4935), .Y(n6362) );
  AOI211X1 U7624 ( .A0(n5092), .A1(n5919), .B0(n6363), .C0(n3350), .Y(n6361)
         );
  OAI222XL U7625 ( .A0(n5921), .A1(n6193), .B0(n5922), .B1(n4980), .C0(n5923), 
        .C1(n4983), .Y(n6363) );
  OAI21XL U7626 ( .A0(n6364), .A1(n5925), .B0(n6365), .Y(n8275) );
  MXI2X1 U7627 ( .A(\ImageBuffer[6][5] ), .B(n4974), .S0(n4936), .Y(n6365) );
  AOI211X1 U7628 ( .A0(n5092), .A1(n5928), .B0(n6366), .C0(n3349), .Y(n6364)
         );
  OAI222XL U7629 ( .A0(n5930), .A1(n4979), .B0(n5931), .B1(n4980), .C0(n5932), 
        .C1(n4983), .Y(n6366) );
  OAI21XL U7630 ( .A0(n6367), .A1(n5934), .B0(n6368), .Y(n8276) );
  MXI2X1 U7631 ( .A(\ImageBuffer[5][5] ), .B(n4976), .S0(n4937), .Y(n6368) );
  AOI211X1 U7632 ( .A0(n5092), .A1(n5937), .B0(n6369), .C0(n6192), .Y(n6367)
         );
  OAI222XL U7633 ( .A0(n5939), .A1(n4978), .B0(n5940), .B1(n4980), .C0(n5941), 
        .C1(n4983), .Y(n6369) );
  OAI21XL U7634 ( .A0(n6370), .A1(n5943), .B0(n6371), .Y(n8277) );
  MXI2X1 U7635 ( .A(\ImageBuffer[4][5] ), .B(n4975), .S0(n4938), .Y(n6371) );
  AOI211X1 U7636 ( .A0(n5092), .A1(n5946), .B0(n6372), .C0(n3350), .Y(n6370)
         );
  OAI222XL U7637 ( .A0(n5948), .A1(n4977), .B0(n5949), .B1(n4980), .C0(n5950), 
        .C1(n4983), .Y(n6372) );
  OAI21XL U7638 ( .A0(n6373), .A1(n5952), .B0(n6374), .Y(n8278) );
  MXI2X1 U7639 ( .A(\ImageBuffer[3][5] ), .B(n4974), .S0(n4939), .Y(n6374) );
  AOI211X1 U7640 ( .A0(n5092), .A1(n5955), .B0(n6375), .C0(n3349), .Y(n6373)
         );
  OAI222XL U7641 ( .A0(n5957), .A1(n4978), .B0(n5958), .B1(n4980), .C0(n5959), 
        .C1(n4983), .Y(n6375) );
  OAI21XL U7642 ( .A0(n6376), .A1(n5961), .B0(n6377), .Y(n8279) );
  MXI2X1 U7643 ( .A(\ImageBuffer[2][5] ), .B(n6190), .S0(n4940), .Y(n6377) );
  AOI211X1 U7644 ( .A0(n5092), .A1(n5964), .B0(n6378), .C0(n3350), .Y(n6376)
         );
  OAI21XL U7645 ( .A0(n6379), .A1(n5970), .B0(n6380), .Y(n8280) );
  MXI2X1 U7646 ( .A(\ImageBuffer[1][5] ), .B(n6190), .S0(n4941), .Y(n6380) );
  AOI211X1 U7647 ( .A0(n5092), .A1(n5973), .B0(n6381), .C0(n6192), .Y(n6379)
         );
  OAI222XL U7648 ( .A0(n5975), .A1(n4979), .B0(n5976), .B1(n4980), .C0(n5977), 
        .C1(n4983), .Y(n6381) );
  MXI2X1 U7649 ( .A(\ImageBuffer[0][5] ), .B(n4976), .S0(n4942), .Y(n6383) );
  NOR2BX1 U7650 ( .AN(IROM_Q[5]), .B(n4945), .Y(n6190) );
  OAI222XL U7651 ( .A0(n5989), .A1(n6193), .B0(n5990), .B1(n4980), .C0(n5991), 
        .C1(n4983), .Y(n6384) );
  CLKINVX1 U7652 ( .A(N2768), .Y(n6194) );
  CLKINVX1 U7653 ( .A(n4869), .Y(n6193) );
  OAI222XL U7654 ( .A0(n5415), .A1(n4991), .B0(n5416), .B1(n4994), .C0(n5418), 
        .C1(n4996), .Y(n6389) );
  OAI222XL U7655 ( .A0(n5426), .A1(n4989), .B0(n5427), .B1(n4994), .C0(n5428), 
        .C1(n4996), .Y(n6396) );
  MXI2X1 U7656 ( .A(\ImageBuffer[61][4] ), .B(n4986), .S0(n4875), .Y(n6398) );
  OAI222XL U7657 ( .A0(n5435), .A1(n4990), .B0(n5436), .B1(n4994), .C0(n5437), 
        .C1(n4995), .Y(n6399) );
  OAI222XL U7658 ( .A0(n5444), .A1(n4989), .B0(n5445), .B1(n4994), .C0(n5446), 
        .C1(n4995), .Y(n6402) );
  OAI222XL U7659 ( .A0(n5453), .A1(n6391), .B0(n5454), .B1(n4993), .C0(n5455), 
        .C1(n4996), .Y(n6405) );
  MXI2X1 U7660 ( .A(\ImageBuffer[58][4] ), .B(n4987), .S0(n4878), .Y(n6407) );
  OAI222XL U7661 ( .A0(n5471), .A1(n6391), .B0(n5472), .B1(n4993), .C0(n5473), 
        .C1(n4995), .Y(n6411) );
  OAI21XL U7662 ( .A0(n6412), .A1(n5475), .B0(n6413), .Y(n8289) );
  AOI211X1 U7663 ( .A0(n5090), .A1(n5478), .B0(n6414), .C0(n3356), .Y(n6412)
         );
  OAI222XL U7664 ( .A0(n5480), .A1(n4989), .B0(n5481), .B1(n4994), .C0(n5482), 
        .C1(n4997), .Y(n6414) );
  OAI222XL U7665 ( .A0(n5489), .A1(n4990), .B0(n5490), .B1(n4994), .C0(n5491), 
        .C1(n4995), .Y(n6417) );
  OAI222XL U7666 ( .A0(n5498), .A1(n6391), .B0(n5499), .B1(n4993), .C0(n5500), 
        .C1(n4996), .Y(n6420) );
  OAI21XL U7667 ( .A0(n6421), .A1(n5502), .B0(n6422), .Y(n8292) );
  AOI211X1 U7668 ( .A0(n5090), .A1(n5505), .B0(n6423), .C0(n3356), .Y(n6421)
         );
  OAI222XL U7669 ( .A0(n5507), .A1(n4989), .B0(n5508), .B1(n4994), .C0(n5509), 
        .C1(n4995), .Y(n6423) );
  OAI21XL U7670 ( .A0(n6424), .A1(n5511), .B0(n6425), .Y(n8293) );
  OAI222XL U7671 ( .A0(n5516), .A1(n4991), .B0(n5517), .B1(n4994), .C0(n5518), 
        .C1(n4996), .Y(n6426) );
  OAI21XL U7672 ( .A0(n6427), .A1(n5520), .B0(n6428), .Y(n8294) );
  OAI222XL U7673 ( .A0(n5525), .A1(n4991), .B0(n5526), .B1(n4992), .C0(n5527), 
        .C1(n4996), .Y(n6429) );
  OAI21XL U7674 ( .A0(n6430), .A1(n5529), .B0(n6431), .Y(n8295) );
  AOI211X1 U7675 ( .A0(n5090), .A1(n5532), .B0(n6432), .C0(n3354), .Y(n6430)
         );
  OAI222XL U7676 ( .A0(n5534), .A1(n6391), .B0(n5535), .B1(n4994), .C0(n5536), 
        .C1(n4996), .Y(n6432) );
  OAI21XL U7677 ( .A0(n6433), .A1(n5538), .B0(n6434), .Y(n8296) );
  OAI222XL U7678 ( .A0(n5543), .A1(n4990), .B0(n5544), .B1(n4993), .C0(n5545), 
        .C1(n4995), .Y(n6435) );
  OAI21XL U7679 ( .A0(n6436), .A1(n5547), .B0(n6437), .Y(n8297) );
  OAI222XL U7680 ( .A0(n5552), .A1(n4989), .B0(n5553), .B1(n4992), .C0(n5554), 
        .C1(n4996), .Y(n6438) );
  OAI21XL U7681 ( .A0(n6439), .A1(n5556), .B0(n6440), .Y(n8298) );
  AOI211X1 U7682 ( .A0(n5090), .A1(n5559), .B0(n6441), .C0(n3355), .Y(n6439)
         );
  OAI222XL U7683 ( .A0(n5561), .A1(n4989), .B0(n5562), .B1(n6392), .C0(n5563), 
        .C1(n4997), .Y(n6441) );
  OAI21XL U7684 ( .A0(n6442), .A1(n5565), .B0(n6443), .Y(n8299) );
  MXI2X1 U7685 ( .A(\ImageBuffer[46][4] ), .B(n4988), .S0(n4892), .Y(n6443) );
  OAI222XL U7686 ( .A0(n5570), .A1(n4989), .B0(n5571), .B1(n4994), .C0(n5572), 
        .C1(n4997), .Y(n6444) );
  OAI21XL U7687 ( .A0(n6445), .A1(n5574), .B0(n6446), .Y(n8300) );
  AOI211X1 U7688 ( .A0(n5090), .A1(n5577), .B0(n6447), .C0(n3354), .Y(n6445)
         );
  OAI222XL U7689 ( .A0(n5579), .A1(n4989), .B0(n5580), .B1(n4993), .C0(n5581), 
        .C1(n4997), .Y(n6447) );
  OAI21XL U7690 ( .A0(n6448), .A1(n5583), .B0(n6449), .Y(n8301) );
  MXI2X1 U7691 ( .A(\ImageBuffer[44][4] ), .B(n4988), .S0(n4894), .Y(n6449) );
  AOI211X1 U7692 ( .A0(n5090), .A1(n5586), .B0(n6450), .C0(n3356), .Y(n6448)
         );
  OAI222XL U7693 ( .A0(n5588), .A1(n4989), .B0(n5589), .B1(n4994), .C0(n5590), 
        .C1(n4997), .Y(n6450) );
  OAI21XL U7694 ( .A0(n6451), .A1(n5592), .B0(n6452), .Y(n8302) );
  AOI211X1 U7695 ( .A0(n5090), .A1(n5595), .B0(n6453), .C0(n3356), .Y(n6451)
         );
  OAI222XL U7696 ( .A0(n5597), .A1(n4989), .B0(n5598), .B1(n6392), .C0(n5599), 
        .C1(n4997), .Y(n6453) );
  OAI21XL U7697 ( .A0(n6454), .A1(n5601), .B0(n6455), .Y(n8303) );
  AOI211X1 U7698 ( .A0(n5090), .A1(n5604), .B0(n6456), .C0(n3355), .Y(n6454)
         );
  OAI222XL U7699 ( .A0(n5606), .A1(n4989), .B0(n5607), .B1(n4994), .C0(n5608), 
        .C1(n4997), .Y(n6456) );
  OAI21XL U7700 ( .A0(n6457), .A1(n5610), .B0(n6458), .Y(n8304) );
  AOI211X1 U7701 ( .A0(n5090), .A1(n5613), .B0(n6459), .C0(n3354), .Y(n6457)
         );
  OAI222XL U7702 ( .A0(n5615), .A1(n4989), .B0(n5616), .B1(n4994), .C0(n5617), 
        .C1(n4997), .Y(n6459) );
  OAI21XL U7703 ( .A0(n6460), .A1(n5619), .B0(n6461), .Y(n8305) );
  OAI222XL U7704 ( .A0(n5624), .A1(n4990), .B0(n5625), .B1(n4994), .C0(n5626), 
        .C1(n4997), .Y(n6462) );
  OAI21XL U7705 ( .A0(n6463), .A1(n5628), .B0(n6464), .Y(n8306) );
  AOI211X1 U7706 ( .A0(n5090), .A1(n5631), .B0(n6465), .C0(n3356), .Y(n6463)
         );
  OAI222XL U7707 ( .A0(n5633), .A1(n4989), .B0(n5634), .B1(n6392), .C0(n5635), 
        .C1(n4997), .Y(n6465) );
  OAI222XL U7708 ( .A0(n5642), .A1(n4991), .B0(n5643), .B1(n4992), .C0(n5644), 
        .C1(n4997), .Y(n6468) );
  OAI21XL U7709 ( .A0(n6469), .A1(n5646), .B0(n6470), .Y(n8308) );
  AOI211X1 U7710 ( .A0(n5090), .A1(n5649), .B0(n6471), .C0(n3355), .Y(n6469)
         );
  OAI222XL U7711 ( .A0(n5651), .A1(n4989), .B0(n5652), .B1(n6392), .C0(n5653), 
        .C1(n4997), .Y(n6471) );
  OAI21XL U7712 ( .A0(n6472), .A1(n5655), .B0(n6473), .Y(n8309) );
  AOI211X1 U7713 ( .A0(n5090), .A1(n5658), .B0(n6474), .C0(n3354), .Y(n6472)
         );
  OAI222XL U7714 ( .A0(n5660), .A1(n4989), .B0(n5661), .B1(n6392), .C0(n5662), 
        .C1(n4997), .Y(n6474) );
  OAI21XL U7715 ( .A0(n6475), .A1(n5664), .B0(n6476), .Y(n8310) );
  OAI222XL U7716 ( .A0(n5669), .A1(n4991), .B0(n5670), .B1(n4993), .C0(n5671), 
        .C1(n4997), .Y(n6477) );
  OAI222XL U7717 ( .A0(n5678), .A1(n4991), .B0(n5679), .B1(n4993), .C0(n5680), 
        .C1(n4997), .Y(n6480) );
  OAI222XL U7718 ( .A0(n5687), .A1(n4991), .B0(n5688), .B1(n4993), .C0(n5689), 
        .C1(n4997), .Y(n6483) );
  OAI21XL U7719 ( .A0(n6484), .A1(n5691), .B0(n6485), .Y(n8313) );
  OAI222XL U7720 ( .A0(n5696), .A1(n4991), .B0(n5697), .B1(n4993), .C0(n5698), 
        .C1(n4997), .Y(n6486) );
  OAI21XL U7721 ( .A0(n6487), .A1(n5700), .B0(n6488), .Y(n8314) );
  OAI222XL U7722 ( .A0(n5705), .A1(n4991), .B0(n5706), .B1(n4993), .C0(n5707), 
        .C1(n4997), .Y(n6489) );
  OAI21XL U7723 ( .A0(n6490), .A1(n5709), .B0(n6491), .Y(n8315) );
  OAI222XL U7724 ( .A0(n5714), .A1(n4991), .B0(n5715), .B1(n4993), .C0(n5716), 
        .C1(n4997), .Y(n6492) );
  OAI21XL U7725 ( .A0(n6493), .A1(n5718), .B0(n6494), .Y(n8316) );
  OAI222XL U7726 ( .A0(n5723), .A1(n4991), .B0(n5724), .B1(n4993), .C0(n5725), 
        .C1(n4997), .Y(n6495) );
  OAI222XL U7727 ( .A0(n5732), .A1(n4991), .B0(n5733), .B1(n4993), .C0(n5734), 
        .C1(n4997), .Y(n6498) );
  OAI21XL U7728 ( .A0(n6499), .A1(n5736), .B0(n6500), .Y(n8318) );
  AOI211X1 U7729 ( .A0(n5090), .A1(n5739), .B0(n6501), .C0(n3355), .Y(n6499)
         );
  OAI222XL U7730 ( .A0(n5741), .A1(n4991), .B0(n5742), .B1(n4993), .C0(n5743), 
        .C1(n4996), .Y(n6501) );
  OAI21XL U7731 ( .A0(n6502), .A1(n5745), .B0(n6503), .Y(n8319) );
  AOI211X1 U7732 ( .A0(n5090), .A1(n5748), .B0(n6504), .C0(n3355), .Y(n6502)
         );
  OAI222XL U7733 ( .A0(n5750), .A1(n4991), .B0(n5751), .B1(n4993), .C0(n5752), 
        .C1(n4995), .Y(n6504) );
  OAI21XL U7734 ( .A0(n6505), .A1(n5754), .B0(n6506), .Y(n8320) );
  AOI211X1 U7735 ( .A0(n5090), .A1(n5757), .B0(n6507), .C0(n3354), .Y(n6505)
         );
  OAI222XL U7736 ( .A0(n5759), .A1(n4991), .B0(n5760), .B1(n4993), .C0(n5761), 
        .C1(n6393), .Y(n6507) );
  OAI21XL U7737 ( .A0(n6508), .A1(n5763), .B0(n6509), .Y(n8321) );
  AOI211X1 U7738 ( .A0(n5090), .A1(n5766), .B0(n6510), .C0(n3356), .Y(n6508)
         );
  OAI222XL U7739 ( .A0(n5768), .A1(n4991), .B0(n5769), .B1(n4993), .C0(n5770), 
        .C1(n4995), .Y(n6510) );
  OAI21XL U7740 ( .A0(n6511), .A1(n5772), .B0(n6512), .Y(n8322) );
  AOI211X1 U7741 ( .A0(n5090), .A1(n5775), .B0(n6513), .C0(n3355), .Y(n6511)
         );
  OAI222XL U7742 ( .A0(n5777), .A1(n4990), .B0(n5778), .B1(n4994), .C0(n5779), 
        .C1(n4996), .Y(n6513) );
  OAI21XL U7743 ( .A0(n6514), .A1(n5781), .B0(n6515), .Y(n8323) );
  AOI211X1 U7744 ( .A0(n5090), .A1(n5784), .B0(n6516), .C0(n3356), .Y(n6514)
         );
  OAI21XL U7745 ( .A0(n6517), .A1(n5790), .B0(n6518), .Y(n8324) );
  AOI211X1 U7746 ( .A0(n5090), .A1(n5793), .B0(n6519), .C0(n3354), .Y(n6517)
         );
  OAI222XL U7747 ( .A0(n5795), .A1(n4989), .B0(n5796), .B1(n4994), .C0(n5797), 
        .C1(n4996), .Y(n6519) );
  OAI21XL U7748 ( .A0(n6520), .A1(n5799), .B0(n6521), .Y(n8325) );
  AOI211X1 U7749 ( .A0(n5090), .A1(n5802), .B0(n6522), .C0(n3355), .Y(n6520)
         );
  OAI222XL U7750 ( .A0(n5804), .A1(n4989), .B0(n5805), .B1(n4994), .C0(n5806), 
        .C1(n4996), .Y(n6522) );
  OAI21XL U7751 ( .A0(n6523), .A1(n5808), .B0(n6524), .Y(n8326) );
  MXI2X1 U7752 ( .A(\ImageBuffer[19][4] ), .B(n4987), .S0(n4922), .Y(n6524) );
  AOI211X1 U7753 ( .A0(n5090), .A1(n5811), .B0(n6525), .C0(n3355), .Y(n6523)
         );
  OAI222XL U7754 ( .A0(n5813), .A1(n4991), .B0(n5814), .B1(n4994), .C0(n5815), 
        .C1(n4996), .Y(n6525) );
  OAI21XL U7755 ( .A0(n6526), .A1(n5817), .B0(n6527), .Y(n8327) );
  AOI211X1 U7756 ( .A0(n5090), .A1(n5820), .B0(n6528), .C0(n3356), .Y(n6526)
         );
  OAI222XL U7757 ( .A0(n5822), .A1(n4989), .B0(n5823), .B1(n4992), .C0(n5824), 
        .C1(n4996), .Y(n6528) );
  OAI222XL U7758 ( .A0(n5831), .A1(n4991), .B0(n5832), .B1(n4994), .C0(n5833), 
        .C1(n4996), .Y(n6531) );
  OAI21XL U7759 ( .A0(n6532), .A1(n5835), .B0(n6533), .Y(n8329) );
  MXI2X1 U7760 ( .A(\ImageBuffer[16][4] ), .B(n4987), .S0(n4925), .Y(n6533) );
  AOI211X1 U7761 ( .A0(n5090), .A1(n5838), .B0(n6534), .C0(n3355), .Y(n6532)
         );
  OAI222XL U7762 ( .A0(n5840), .A1(n4991), .B0(n5841), .B1(n4992), .C0(n5842), 
        .C1(n4996), .Y(n6534) );
  OAI21XL U7763 ( .A0(n6535), .A1(n5844), .B0(n6536), .Y(n8330) );
  AOI211X1 U7764 ( .A0(n5090), .A1(n5847), .B0(n6537), .C0(n3355), .Y(n6535)
         );
  OAI222XL U7765 ( .A0(n5849), .A1(n4991), .B0(n5850), .B1(n4992), .C0(n5851), 
        .C1(n4996), .Y(n6537) );
  OAI21XL U7766 ( .A0(n6538), .A1(n5853), .B0(n6539), .Y(n8331) );
  AOI211X1 U7767 ( .A0(n5090), .A1(n5856), .B0(n6540), .C0(n3356), .Y(n6538)
         );
  OAI222XL U7768 ( .A0(n5858), .A1(n4990), .B0(n5859), .B1(n4994), .C0(n5860), 
        .C1(n4996), .Y(n6540) );
  OAI21XL U7769 ( .A0(n6541), .A1(n5862), .B0(n6542), .Y(n8332) );
  AOI211X1 U7770 ( .A0(n5090), .A1(n5865), .B0(n6543), .C0(n3354), .Y(n6541)
         );
  OAI222XL U7771 ( .A0(n5867), .A1(n4990), .B0(n5868), .B1(n4992), .C0(n5869), 
        .C1(n4996), .Y(n6543) );
  OAI21XL U7772 ( .A0(n6544), .A1(n5871), .B0(n6545), .Y(n8333) );
  AOI211X1 U7773 ( .A0(n5090), .A1(n5874), .B0(n6546), .C0(n3355), .Y(n6544)
         );
  OAI222XL U7774 ( .A0(n5876), .A1(n6391), .B0(n5877), .B1(n4992), .C0(n5878), 
        .C1(n4996), .Y(n6546) );
  OAI21XL U7775 ( .A0(n6547), .A1(n5880), .B0(n6548), .Y(n8334) );
  MXI2X1 U7776 ( .A(\ImageBuffer[11][4] ), .B(n4986), .S0(n4931), .Y(n6548) );
  AOI211X1 U7777 ( .A0(n5090), .A1(n5883), .B0(n6549), .C0(n3354), .Y(n6547)
         );
  OAI222XL U7778 ( .A0(n5885), .A1(n4990), .B0(n5886), .B1(n4992), .C0(n5887), 
        .C1(n4995), .Y(n6549) );
  OAI21XL U7779 ( .A0(n6550), .A1(n5889), .B0(n6551), .Y(n8335) );
  MXI2X1 U7780 ( .A(\ImageBuffer[10][4] ), .B(n4986), .S0(n4932), .Y(n6551) );
  AOI211X1 U7781 ( .A0(n5090), .A1(n5892), .B0(n6552), .C0(n3356), .Y(n6550)
         );
  OAI222XL U7782 ( .A0(n5894), .A1(n4990), .B0(n5895), .B1(n4992), .C0(n5896), 
        .C1(n4995), .Y(n6552) );
  OAI21XL U7783 ( .A0(n6553), .A1(n5898), .B0(n6554), .Y(n8336) );
  MXI2X1 U7784 ( .A(\ImageBuffer[9][4] ), .B(n4986), .S0(n4933), .Y(n6554) );
  AOI211X1 U7785 ( .A0(n5090), .A1(n5901), .B0(n6555), .C0(n3355), .Y(n6553)
         );
  OAI222XL U7786 ( .A0(n5903), .A1(n4990), .B0(n5904), .B1(n4992), .C0(n5905), 
        .C1(n4995), .Y(n6555) );
  OAI21XL U7787 ( .A0(n6556), .A1(n5907), .B0(n6557), .Y(n8337) );
  MXI2X1 U7788 ( .A(\ImageBuffer[8][4] ), .B(n4986), .S0(n4934), .Y(n6557) );
  AOI211X1 U7789 ( .A0(n5090), .A1(n5910), .B0(n6558), .C0(n3354), .Y(n6556)
         );
  OAI222XL U7790 ( .A0(n5912), .A1(n4990), .B0(n5913), .B1(n4992), .C0(n5914), 
        .C1(n4995), .Y(n6558) );
  OAI21XL U7791 ( .A0(n6559), .A1(n5916), .B0(n6560), .Y(n8338) );
  MXI2X1 U7792 ( .A(\ImageBuffer[7][4] ), .B(n4986), .S0(n4935), .Y(n6560) );
  AOI211X1 U7793 ( .A0(n5090), .A1(n5919), .B0(n6561), .C0(n3356), .Y(n6559)
         );
  OAI222XL U7794 ( .A0(n5921), .A1(n4990), .B0(n5922), .B1(n4992), .C0(n5923), 
        .C1(n4995), .Y(n6561) );
  OAI21XL U7795 ( .A0(n6562), .A1(n5925), .B0(n6563), .Y(n8339) );
  MXI2X1 U7796 ( .A(\ImageBuffer[6][4] ), .B(n4986), .S0(n4936), .Y(n6563) );
  AOI211X1 U7797 ( .A0(n5090), .A1(n5928), .B0(n6564), .C0(n3355), .Y(n6562)
         );
  OAI222XL U7798 ( .A0(n5930), .A1(n4990), .B0(n5931), .B1(n4992), .C0(n5932), 
        .C1(n4995), .Y(n6564) );
  OAI21XL U7799 ( .A0(n6565), .A1(n5934), .B0(n6566), .Y(n8340) );
  MXI2X1 U7800 ( .A(\ImageBuffer[5][4] ), .B(n4986), .S0(n4937), .Y(n6566) );
  AOI211X1 U7801 ( .A0(n5090), .A1(n5937), .B0(n6567), .C0(n3354), .Y(n6565)
         );
  OAI222XL U7802 ( .A0(n5939), .A1(n4990), .B0(n5940), .B1(n4992), .C0(n5941), 
        .C1(n4995), .Y(n6567) );
  OAI21XL U7803 ( .A0(n6568), .A1(n5943), .B0(n6569), .Y(n8341) );
  MXI2X1 U7804 ( .A(\ImageBuffer[4][4] ), .B(n4986), .S0(n4938), .Y(n6569) );
  AOI211X1 U7805 ( .A0(n5090), .A1(n5946), .B0(n6570), .C0(n3356), .Y(n6568)
         );
  OAI222XL U7806 ( .A0(n5948), .A1(n4990), .B0(n5949), .B1(n4992), .C0(n5950), 
        .C1(n4995), .Y(n6570) );
  OAI21XL U7807 ( .A0(n6571), .A1(n5952), .B0(n6572), .Y(n8342) );
  MXI2X1 U7808 ( .A(\ImageBuffer[3][4] ), .B(n4986), .S0(n4939), .Y(n6572) );
  AOI211X1 U7809 ( .A0(n5090), .A1(n5955), .B0(n6573), .C0(n3355), .Y(n6571)
         );
  OAI222XL U7810 ( .A0(n5957), .A1(n4990), .B0(n5958), .B1(n4992), .C0(n5959), 
        .C1(n4995), .Y(n6573) );
  OAI21XL U7811 ( .A0(n6574), .A1(n5961), .B0(n6575), .Y(n8343) );
  MXI2X1 U7812 ( .A(\ImageBuffer[2][4] ), .B(n4986), .S0(n4940), .Y(n6575) );
  AOI211X1 U7813 ( .A0(n5090), .A1(n5964), .B0(n6576), .C0(n3354), .Y(n6574)
         );
  OAI21XL U7814 ( .A0(n6577), .A1(n5970), .B0(n6578), .Y(n8344) );
  MXI2X1 U7815 ( .A(\ImageBuffer[1][4] ), .B(n4986), .S0(n4941), .Y(n6578) );
  AOI211X1 U7816 ( .A0(n5090), .A1(n5973), .B0(n6579), .C0(n3354), .Y(n6577)
         );
  OAI222XL U7817 ( .A0(n5975), .A1(n4990), .B0(n5976), .B1(n4992), .C0(n5977), 
        .C1(n4995), .Y(n6579) );
  MXI2X1 U7818 ( .A(\ImageBuffer[0][4] ), .B(n4986), .S0(n4942), .Y(n6581) );
  NOR2BX1 U7819 ( .AN(IROM_Q[4]), .B(n4945), .Y(n6388) );
  OAI222XL U7820 ( .A0(n5989), .A1(n4990), .B0(n5990), .B1(n4992), .C0(n5991), 
        .C1(n4995), .Y(n6582) );
  CLKINVX1 U7821 ( .A(N2769), .Y(n6392) );
  CLKINVX1 U7822 ( .A(n4870), .Y(n6391) );
  OAI222XL U7823 ( .A0(n5415), .A1(n5004), .B0(n5416), .B1(n5006), .C0(n5418), 
        .C1(n5010), .Y(n6587) );
  OAI222XL U7824 ( .A0(n5426), .A1(n5003), .B0(n5427), .B1(n5005), .C0(n5428), 
        .C1(n5008), .Y(n6593) );
  OAI222XL U7825 ( .A0(n5435), .A1(n5003), .B0(n5436), .B1(n5007), .C0(n5437), 
        .C1(n5008), .Y(n6596) );
  OAI222XL U7826 ( .A0(n5444), .A1(n5002), .B0(n5445), .B1(n5005), .C0(n5446), 
        .C1(n5008), .Y(n6599) );
  MXI2X1 U7827 ( .A(\ImageBuffer[59][3] ), .B(n5001), .S0(n4877), .Y(n6601) );
  OAI222XL U7828 ( .A0(n5453), .A1(n5004), .B0(n5454), .B1(n5005), .C0(n5455), 
        .C1(n5010), .Y(n6602) );
  MXI2X1 U7829 ( .A(\ImageBuffer[58][3] ), .B(n5001), .S0(n4878), .Y(n6604) );
  OAI222XL U7830 ( .A0(n5462), .A1(n5003), .B0(n5463), .B1(n5006), .C0(n5464), 
        .C1(n5010), .Y(n6605) );
  MXI2X1 U7831 ( .A(\ImageBuffer[57][3] ), .B(n5001), .S0(n4879), .Y(n6607) );
  OAI222XL U7832 ( .A0(n5471), .A1(n5003), .B0(n5472), .B1(n5007), .C0(n5473), 
        .C1(n5010), .Y(n6608) );
  MXI2X1 U7833 ( .A(\ImageBuffer[56][3] ), .B(n5001), .S0(n4880), .Y(n6610) );
  OAI222XL U7834 ( .A0(n5480), .A1(n5002), .B0(n5481), .B1(n6590), .C0(n5482), 
        .C1(n5010), .Y(n6611) );
  MXI2X1 U7835 ( .A(\ImageBuffer[55][3] ), .B(n5001), .S0(n4882), .Y(n6613) );
  OAI222XL U7836 ( .A0(n5489), .A1(n5003), .B0(n5490), .B1(n6590), .C0(n5491), 
        .C1(n5010), .Y(n6614) );
  MXI2X1 U7837 ( .A(\ImageBuffer[54][3] ), .B(n5001), .S0(n4883), .Y(n6616) );
  MXI2X1 U7838 ( .A(\ImageBuffer[53][3] ), .B(n5001), .S0(n4884), .Y(n6619) );
  OAI222XL U7839 ( .A0(n5507), .A1(n5004), .B0(n5508), .B1(n6590), .C0(n5509), 
        .C1(n5010), .Y(n6620) );
  MXI2X1 U7840 ( .A(\ImageBuffer[52][3] ), .B(n5001), .S0(n4885), .Y(n6622) );
  OAI222XL U7841 ( .A0(n5516), .A1(n5003), .B0(n5517), .B1(n5007), .C0(n5518), 
        .C1(n5010), .Y(n6623) );
  MXI2X1 U7842 ( .A(\ImageBuffer[51][3] ), .B(n5001), .S0(n4886), .Y(n6625) );
  OAI222XL U7843 ( .A0(n5525), .A1(n5002), .B0(n5526), .B1(n5007), .C0(n5527), 
        .C1(n5010), .Y(n6626) );
  MXI2X1 U7844 ( .A(\ImageBuffer[50][3] ), .B(n5001), .S0(n4887), .Y(n6628) );
  OAI222XL U7845 ( .A0(n5534), .A1(n5003), .B0(n5535), .B1(n5005), .C0(n5536), 
        .C1(n5010), .Y(n6629) );
  MXI2X1 U7846 ( .A(\ImageBuffer[49][3] ), .B(n5001), .S0(n4888), .Y(n6631) );
  OAI222XL U7847 ( .A0(n5543), .A1(n5004), .B0(n5544), .B1(n5006), .C0(n5545), 
        .C1(n5010), .Y(n6632) );
  MXI2X1 U7848 ( .A(\ImageBuffer[48][3] ), .B(n5001), .S0(n4889), .Y(n6634) );
  OAI222XL U7849 ( .A0(n5552), .A1(n5002), .B0(n5553), .B1(n5006), .C0(n5554), 
        .C1(n5010), .Y(n6635) );
  MXI2X1 U7850 ( .A(\ImageBuffer[47][3] ), .B(n5000), .S0(n4891), .Y(n6637) );
  OAI222XL U7851 ( .A0(n5561), .A1(n5003), .B0(n5562), .B1(n5007), .C0(n5563), 
        .C1(n5009), .Y(n6638) );
  MXI2X1 U7852 ( .A(\ImageBuffer[46][3] ), .B(n5000), .S0(n4892), .Y(n6640) );
  OAI222XL U7853 ( .A0(n5570), .A1(n5004), .B0(n5571), .B1(n5007), .C0(n5572), 
        .C1(n5008), .Y(n6641) );
  MXI2X1 U7854 ( .A(\ImageBuffer[45][3] ), .B(n5000), .S0(n4893), .Y(n6643) );
  AOI211X1 U7855 ( .A0(n5084), .A1(n5577), .B0(n6644), .C0(n6588), .Y(n6642)
         );
  OAI222XL U7856 ( .A0(n5579), .A1(n5002), .B0(n5580), .B1(n5007), .C0(n5581), 
        .C1(n5008), .Y(n6644) );
  MXI2X1 U7857 ( .A(\ImageBuffer[44][3] ), .B(n5000), .S0(n4894), .Y(n6646) );
  OAI222XL U7858 ( .A0(n5588), .A1(n5003), .B0(n5589), .B1(n5007), .C0(n5590), 
        .C1(n5010), .Y(n6647) );
  MXI2X1 U7859 ( .A(\ImageBuffer[43][3] ), .B(n5000), .S0(n4895), .Y(n6649) );
  OAI222XL U7860 ( .A0(n5597), .A1(n5004), .B0(n5598), .B1(n5007), .C0(n5599), 
        .C1(n5009), .Y(n6650) );
  MXI2X1 U7861 ( .A(\ImageBuffer[42][3] ), .B(n5000), .S0(n4896), .Y(n6652) );
  OAI222XL U7862 ( .A0(n5606), .A1(n5002), .B0(n5607), .B1(n5007), .C0(n5608), 
        .C1(n5010), .Y(n6653) );
  MXI2X1 U7863 ( .A(\ImageBuffer[41][3] ), .B(n5000), .S0(n4897), .Y(n6655) );
  OAI222XL U7864 ( .A0(n5615), .A1(n5003), .B0(n5616), .B1(n5007), .C0(n5617), 
        .C1(n5010), .Y(n6656) );
  MXI2X1 U7865 ( .A(\ImageBuffer[40][3] ), .B(n5000), .S0(n4898), .Y(n6658) );
  OAI222XL U7866 ( .A0(n5624), .A1(n5004), .B0(n5625), .B1(n5007), .C0(n5626), 
        .C1(n5008), .Y(n6659) );
  MXI2X1 U7867 ( .A(\ImageBuffer[39][3] ), .B(n5000), .S0(n4900), .Y(n6661) );
  OAI222XL U7868 ( .A0(n5633), .A1(n5002), .B0(n5634), .B1(n5007), .C0(n5635), 
        .C1(n5010), .Y(n6662) );
  MXI2X1 U7869 ( .A(\ImageBuffer[38][3] ), .B(n5000), .S0(n4901), .Y(n6664) );
  OAI222XL U7870 ( .A0(n5642), .A1(n5003), .B0(n5643), .B1(n5007), .C0(n5644), 
        .C1(n5010), .Y(n6665) );
  MXI2X1 U7871 ( .A(\ImageBuffer[37][3] ), .B(n5000), .S0(n4902), .Y(n6667) );
  OAI222XL U7872 ( .A0(n5651), .A1(n5004), .B0(n5652), .B1(n5007), .C0(n5653), 
        .C1(n5008), .Y(n6668) );
  MXI2X1 U7873 ( .A(\ImageBuffer[36][3] ), .B(n5000), .S0(n4903), .Y(n6670) );
  OAI222XL U7874 ( .A0(n5660), .A1(n5002), .B0(n5661), .B1(n5007), .C0(n5662), 
        .C1(n5008), .Y(n6671) );
  MXI2X1 U7875 ( .A(\ImageBuffer[35][3] ), .B(n4999), .S0(n4904), .Y(n6673) );
  AOI211X1 U7876 ( .A0(n5084), .A1(n5667), .B0(n6674), .C0(n6588), .Y(n6672)
         );
  OAI222XL U7877 ( .A0(n5669), .A1(n5003), .B0(n5670), .B1(n5007), .C0(n5671), 
        .C1(n5009), .Y(n6674) );
  MXI2X1 U7878 ( .A(\ImageBuffer[34][3] ), .B(n4999), .S0(n4905), .Y(n6676) );
  OAI222XL U7879 ( .A0(n5678), .A1(n5004), .B0(n5679), .B1(n5006), .C0(n5680), 
        .C1(n5009), .Y(n6677) );
  MXI2X1 U7880 ( .A(\ImageBuffer[33][3] ), .B(n4999), .S0(n4906), .Y(n6679) );
  AOI211X1 U7881 ( .A0(n5084), .A1(n5685), .B0(n6680), .C0(n3359), .Y(n6678)
         );
  OAI222XL U7882 ( .A0(n5687), .A1(n5004), .B0(n5688), .B1(n5005), .C0(n5689), 
        .C1(n5009), .Y(n6680) );
  MXI2X1 U7883 ( .A(\ImageBuffer[32][3] ), .B(n4999), .S0(n4907), .Y(n6682) );
  OAI222XL U7884 ( .A0(n5696), .A1(n5004), .B0(n5697), .B1(n5007), .C0(n5698), 
        .C1(n5009), .Y(n6683) );
  MXI2X1 U7885 ( .A(\ImageBuffer[31][3] ), .B(n4999), .S0(n4909), .Y(n6685) );
  OAI222XL U7886 ( .A0(n5705), .A1(n5002), .B0(n5706), .B1(n6590), .C0(n5707), 
        .C1(n5009), .Y(n6686) );
  MXI2X1 U7887 ( .A(\ImageBuffer[30][3] ), .B(n4999), .S0(n4910), .Y(n6688) );
  OAI222XL U7888 ( .A0(n5714), .A1(n5002), .B0(n5715), .B1(n5005), .C0(n5716), 
        .C1(n5009), .Y(n6689) );
  MXI2X1 U7889 ( .A(\ImageBuffer[29][3] ), .B(n4999), .S0(n4911), .Y(n6691) );
  OAI222XL U7890 ( .A0(n5723), .A1(n5002), .B0(n5724), .B1(n5007), .C0(n5725), 
        .C1(n5009), .Y(n6692) );
  MXI2X1 U7891 ( .A(\ImageBuffer[28][3] ), .B(n4999), .S0(n4912), .Y(n6694) );
  OAI222XL U7892 ( .A0(n5732), .A1(n5004), .B0(n5733), .B1(n5005), .C0(n5734), 
        .C1(n5009), .Y(n6695) );
  MXI2X1 U7893 ( .A(\ImageBuffer[27][3] ), .B(n4999), .S0(n4913), .Y(n6697) );
  OAI222XL U7894 ( .A0(n5741), .A1(n5004), .B0(n5742), .B1(n5006), .C0(n5743), 
        .C1(n5009), .Y(n6698) );
  MXI2X1 U7895 ( .A(\ImageBuffer[26][3] ), .B(n4999), .S0(n4914), .Y(n6700) );
  OAI222XL U7896 ( .A0(n5750), .A1(n5002), .B0(n5751), .B1(n5005), .C0(n5752), 
        .C1(n5009), .Y(n6701) );
  MXI2X1 U7897 ( .A(\ImageBuffer[25][3] ), .B(n4999), .S0(n4915), .Y(n6703) );
  OAI222XL U7898 ( .A0(n5759), .A1(n5003), .B0(n5760), .B1(n5006), .C0(n5761), 
        .C1(n5009), .Y(n6704) );
  MXI2X1 U7899 ( .A(\ImageBuffer[24][3] ), .B(n4999), .S0(n4916), .Y(n6706) );
  OAI222XL U7900 ( .A0(n5768), .A1(n5003), .B0(n5769), .B1(n5007), .C0(n5770), 
        .C1(n5009), .Y(n6707) );
  MXI2X1 U7901 ( .A(\ImageBuffer[23][3] ), .B(n5001), .S0(n4918), .Y(n6709) );
  OAI222XL U7902 ( .A0(n5777), .A1(n5004), .B0(n5778), .B1(n5006), .C0(n5779), 
        .C1(n5008), .Y(n6710) );
  MXI2X1 U7903 ( .A(\ImageBuffer[22][3] ), .B(n4999), .S0(n4919), .Y(n6712) );
  OAI222XL U7904 ( .A0(n5786), .A1(n5002), .B0(n5787), .B1(n5006), .C0(n5788), 
        .C1(n5008), .Y(n6713) );
  MXI2X1 U7905 ( .A(\ImageBuffer[21][3] ), .B(n5001), .S0(n4920), .Y(n6715) );
  OAI222XL U7906 ( .A0(n5795), .A1(n5003), .B0(n5796), .B1(n5006), .C0(n5797), 
        .C1(n5008), .Y(n6716) );
  MXI2X1 U7907 ( .A(\ImageBuffer[20][3] ), .B(n5001), .S0(n4921), .Y(n6718) );
  OAI222XL U7908 ( .A0(n5804), .A1(n5004), .B0(n5805), .B1(n5006), .C0(n5806), 
        .C1(n5008), .Y(n6719) );
  MXI2X1 U7909 ( .A(\ImageBuffer[19][3] ), .B(n5001), .S0(n4922), .Y(n6721) );
  OAI222XL U7910 ( .A0(n5813), .A1(n5002), .B0(n5814), .B1(n5006), .C0(n5815), 
        .C1(n5008), .Y(n6722) );
  MXI2X1 U7911 ( .A(\ImageBuffer[18][3] ), .B(n4999), .S0(n4923), .Y(n6724) );
  OAI222XL U7912 ( .A0(n5822), .A1(n5003), .B0(n5823), .B1(n5006), .C0(n5824), 
        .C1(n5008), .Y(n6725) );
  MXI2X1 U7913 ( .A(\ImageBuffer[17][3] ), .B(n5001), .S0(n4924), .Y(n6727) );
  OAI222XL U7914 ( .A0(n5831), .A1(n5004), .B0(n5832), .B1(n5006), .C0(n5833), 
        .C1(n5008), .Y(n6728) );
  MXI2X1 U7915 ( .A(\ImageBuffer[16][3] ), .B(n4999), .S0(n4925), .Y(n6730) );
  OAI222XL U7916 ( .A0(n5840), .A1(n5002), .B0(n5841), .B1(n5006), .C0(n5842), 
        .C1(n5008), .Y(n6731) );
  MXI2X1 U7917 ( .A(\ImageBuffer[15][3] ), .B(n4999), .S0(n4927), .Y(n6733) );
  OAI222XL U7918 ( .A0(n5849), .A1(n5003), .B0(n5850), .B1(n5006), .C0(n5851), 
        .C1(n5008), .Y(n6734) );
  MXI2X1 U7919 ( .A(\ImageBuffer[14][3] ), .B(n5001), .S0(n4928), .Y(n6736) );
  OAI222XL U7920 ( .A0(n5858), .A1(n5004), .B0(n5859), .B1(n5006), .C0(n5860), 
        .C1(n5008), .Y(n6737) );
  MXI2X1 U7921 ( .A(\ImageBuffer[13][3] ), .B(n4999), .S0(n4929), .Y(n6739) );
  OAI222XL U7922 ( .A0(n5867), .A1(n5002), .B0(n5868), .B1(n5006), .C0(n5869), 
        .C1(n5008), .Y(n6740) );
  MXI2X1 U7923 ( .A(\ImageBuffer[12][3] ), .B(n4999), .S0(n4930), .Y(n6742) );
  OAI222XL U7924 ( .A0(n5876), .A1(n5003), .B0(n5877), .B1(n5006), .C0(n5878), 
        .C1(n5008), .Y(n6743) );
  MXI2X1 U7925 ( .A(\ImageBuffer[11][3] ), .B(n4998), .S0(n4931), .Y(n6745) );
  OAI222XL U7926 ( .A0(n5885), .A1(n5002), .B0(n5886), .B1(n5005), .C0(n5887), 
        .C1(n5009), .Y(n6746) );
  MXI2X1 U7927 ( .A(\ImageBuffer[10][3] ), .B(n4998), .S0(n4932), .Y(n6748) );
  OAI222XL U7928 ( .A0(n5894), .A1(n5003), .B0(n5895), .B1(n5005), .C0(n5896), 
        .C1(n5009), .Y(n6749) );
  MXI2X1 U7929 ( .A(\ImageBuffer[9][3] ), .B(n4998), .S0(n4933), .Y(n6751) );
  OAI222XL U7930 ( .A0(n5903), .A1(n5004), .B0(n5904), .B1(n5005), .C0(n5905), 
        .C1(n5009), .Y(n6752) );
  MXI2X1 U7931 ( .A(\ImageBuffer[8][3] ), .B(n4998), .S0(n4934), .Y(n6754) );
  OAI222XL U7932 ( .A0(n5912), .A1(n5002), .B0(n5913), .B1(n5005), .C0(n5914), 
        .C1(n5009), .Y(n6755) );
  MXI2X1 U7933 ( .A(\ImageBuffer[7][3] ), .B(n4998), .S0(n4935), .Y(n6757) );
  OAI222XL U7934 ( .A0(n5921), .A1(n5003), .B0(n5922), .B1(n5005), .C0(n5923), 
        .C1(n5009), .Y(n6758) );
  MXI2X1 U7935 ( .A(\ImageBuffer[6][3] ), .B(n4998), .S0(n4936), .Y(n6760) );
  OAI222XL U7936 ( .A0(n5930), .A1(n5004), .B0(n5931), .B1(n5005), .C0(n5932), 
        .C1(n5008), .Y(n6761) );
  MXI2X1 U7937 ( .A(\ImageBuffer[5][3] ), .B(n4998), .S0(n4937), .Y(n6763) );
  OAI222XL U7938 ( .A0(n5939), .A1(n5002), .B0(n5940), .B1(n5005), .C0(n5941), 
        .C1(n5009), .Y(n6764) );
  MXI2X1 U7939 ( .A(\ImageBuffer[4][3] ), .B(n4998), .S0(n4938), .Y(n6766) );
  OAI222XL U7940 ( .A0(n5948), .A1(n5003), .B0(n5949), .B1(n5005), .C0(n5950), 
        .C1(n5010), .Y(n6767) );
  MXI2X1 U7941 ( .A(\ImageBuffer[3][3] ), .B(n4998), .S0(n4939), .Y(n6769) );
  OAI222XL U7942 ( .A0(n5957), .A1(n5004), .B0(n5958), .B1(n5005), .C0(n5959), 
        .C1(n5010), .Y(n6770) );
  MXI2X1 U7943 ( .A(\ImageBuffer[2][3] ), .B(n4998), .S0(n4940), .Y(n6772) );
  MXI2X1 U7944 ( .A(\ImageBuffer[1][3] ), .B(n4998), .S0(n4941), .Y(n6775) );
  OAI222XL U7945 ( .A0(n5975), .A1(n5002), .B0(n5976), .B1(n5005), .C0(n5977), 
        .C1(n5009), .Y(n6776) );
  MXI2X1 U7946 ( .A(\ImageBuffer[0][3] ), .B(n4998), .S0(n4942), .Y(n6778) );
  NOR2BX1 U7947 ( .AN(IROM_Q[3]), .B(n4945), .Y(n6586) );
  AOI211X1 U7948 ( .A0(n5084), .A1(n5983), .B0(n6779), .C0(n3359), .Y(n6777)
         );
  OAI222XL U7949 ( .A0(n5989), .A1(n5002), .B0(n5990), .B1(n5005), .C0(n5991), 
        .C1(n5218), .Y(n6779) );
  CLKINVX1 U7950 ( .A(N2770), .Y(n6590) );
  OAI21XL U7951 ( .A0(n6781), .A1(n5408), .B0(n6782), .Y(n8410) );
  MXI2X1 U7952 ( .A(\ImageBuffer[63][2] ), .B(n5012), .S0(n5411), .Y(n6782) );
  AOI211X1 U7953 ( .A0(n5082), .A1(n5412), .B0(n6784), .C0(n6785), .Y(n6781)
         );
  OAI222XL U7954 ( .A0(n5415), .A1(n5017), .B0(n5416), .B1(n5019), .C0(n5418), 
        .C1(n5021), .Y(n6784) );
  OAI21XL U7955 ( .A0(n6788), .A1(n5421), .B0(n6789), .Y(n8411) );
  MXI2X1 U7956 ( .A(\ImageBuffer[62][2] ), .B(n5011), .S0(n4874), .Y(n6789) );
  AOI211X1 U7957 ( .A0(n5082), .A1(n5424), .B0(n6790), .C0(n6785), .Y(n6788)
         );
  OAI222XL U7958 ( .A0(n5426), .A1(n5016), .B0(n5427), .B1(n5019), .C0(n5428), 
        .C1(n5022), .Y(n6790) );
  MXI2X1 U7959 ( .A(\ImageBuffer[61][2] ), .B(n5011), .S0(n4875), .Y(n6792) );
  AOI211X1 U7960 ( .A0(n5082), .A1(n5433), .B0(n6793), .C0(n6785), .Y(n6791)
         );
  OAI222XL U7961 ( .A0(n5435), .A1(n5015), .B0(n5436), .B1(n5019), .C0(n5437), 
        .C1(n5021), .Y(n6793) );
  OAI21XL U7962 ( .A0(n6794), .A1(n5439), .B0(n6795), .Y(n8413) );
  MXI2X1 U7963 ( .A(\ImageBuffer[60][2] ), .B(n5012), .S0(n4876), .Y(n6795) );
  AOI211X1 U7964 ( .A0(n5082), .A1(n5442), .B0(n6796), .C0(n6785), .Y(n6794)
         );
  OAI222XL U7965 ( .A0(n5444), .A1(n5017), .B0(n5445), .B1(n5018), .C0(n5446), 
        .C1(n5021), .Y(n6796) );
  OAI21XL U7966 ( .A0(n6797), .A1(n5448), .B0(n6798), .Y(n8414) );
  MXI2X1 U7967 ( .A(\ImageBuffer[59][2] ), .B(n5014), .S0(n4877), .Y(n6798) );
  AOI211X1 U7968 ( .A0(n5082), .A1(n5451), .B0(n6799), .C0(n6785), .Y(n6797)
         );
  OAI222XL U7969 ( .A0(n5453), .A1(n5017), .B0(n5454), .B1(n5020), .C0(n5455), 
        .C1(n5024), .Y(n6799) );
  OAI21XL U7970 ( .A0(n6800), .A1(n5457), .B0(n6801), .Y(n8415) );
  MXI2X1 U7971 ( .A(\ImageBuffer[58][2] ), .B(n5014), .S0(n4878), .Y(n6801) );
  AOI211X1 U7972 ( .A0(n5082), .A1(n5460), .B0(n6802), .C0(n6785), .Y(n6800)
         );
  OAI222XL U7973 ( .A0(n5462), .A1(n5017), .B0(n5463), .B1(n5018), .C0(n5464), 
        .C1(n5024), .Y(n6802) );
  OAI21XL U7974 ( .A0(n6803), .A1(n5466), .B0(n6804), .Y(n8416) );
  MXI2X1 U7975 ( .A(\ImageBuffer[57][2] ), .B(n5014), .S0(n4879), .Y(n6804) );
  AOI211X1 U7976 ( .A0(n5082), .A1(n5469), .B0(n6805), .C0(n6785), .Y(n6803)
         );
  OAI222XL U7977 ( .A0(n5471), .A1(n5017), .B0(n5472), .B1(n6787), .C0(n5473), 
        .C1(n5024), .Y(n6805) );
  MXI2X1 U7978 ( .A(\ImageBuffer[56][2] ), .B(n5014), .S0(n4880), .Y(n6807) );
  AOI211X1 U7979 ( .A0(n5082), .A1(n5478), .B0(n6808), .C0(n6785), .Y(n6806)
         );
  MXI2X1 U7980 ( .A(\ImageBuffer[55][2] ), .B(n5014), .S0(n4882), .Y(n6810) );
  MXI2X1 U7981 ( .A(\ImageBuffer[54][2] ), .B(n5014), .S0(n4883), .Y(n6813) );
  OAI222XL U7982 ( .A0(n5498), .A1(n5017), .B0(n5499), .B1(n5020), .C0(n5500), 
        .C1(n5024), .Y(n6814) );
  MXI2X1 U7983 ( .A(\ImageBuffer[53][2] ), .B(n5014), .S0(n4884), .Y(n6816) );
  MXI2X1 U7984 ( .A(\ImageBuffer[52][2] ), .B(n5014), .S0(n4885), .Y(n6819) );
  OAI222XL U7985 ( .A0(n5516), .A1(n5017), .B0(n5517), .B1(n5018), .C0(n5518), 
        .C1(n5024), .Y(n6820) );
  MXI2X1 U7986 ( .A(\ImageBuffer[51][2] ), .B(n5014), .S0(n4886), .Y(n6822) );
  OAI222XL U7987 ( .A0(n5525), .A1(n5017), .B0(n5526), .B1(n6787), .C0(n5527), 
        .C1(n5024), .Y(n6823) );
  MXI2X1 U7988 ( .A(\ImageBuffer[50][2] ), .B(n5014), .S0(n4887), .Y(n6825) );
  MXI2X1 U7989 ( .A(\ImageBuffer[49][2] ), .B(n5014), .S0(n4888), .Y(n6828) );
  OAI222XL U7990 ( .A0(n5543), .A1(n5017), .B0(n5544), .B1(n5019), .C0(n5545), 
        .C1(n5024), .Y(n6829) );
  MXI2X1 U7991 ( .A(\ImageBuffer[48][2] ), .B(n5014), .S0(n4889), .Y(n6831) );
  OAI222XL U7992 ( .A0(n5552), .A1(n5017), .B0(n5553), .B1(n5018), .C0(n5554), 
        .C1(n5024), .Y(n6832) );
  MXI2X1 U7993 ( .A(\ImageBuffer[47][2] ), .B(n5013), .S0(n4891), .Y(n6834) );
  OAI222XL U7994 ( .A0(n5561), .A1(n5016), .B0(n5562), .B1(n5020), .C0(n5563), 
        .C1(n5022), .Y(n6835) );
  MXI2X1 U7995 ( .A(\ImageBuffer[46][2] ), .B(n5013), .S0(n4892), .Y(n6837) );
  OAI222XL U7996 ( .A0(n5570), .A1(n5016), .B0(n5571), .B1(n5020), .C0(n5572), 
        .C1(n5021), .Y(n6838) );
  MXI2X1 U7997 ( .A(\ImageBuffer[45][2] ), .B(n5013), .S0(n4893), .Y(n6840) );
  OAI222XL U7998 ( .A0(n5579), .A1(n5016), .B0(n5580), .B1(n5020), .C0(n5581), 
        .C1(n5023), .Y(n6841) );
  MXI2X1 U7999 ( .A(\ImageBuffer[44][2] ), .B(n5013), .S0(n4894), .Y(n6843) );
  OAI222XL U8000 ( .A0(n5588), .A1(n5016), .B0(n5589), .B1(n5020), .C0(n5590), 
        .C1(n5021), .Y(n6844) );
  MXI2X1 U8001 ( .A(\ImageBuffer[43][2] ), .B(n5013), .S0(n4895), .Y(n6846) );
  OAI222XL U8002 ( .A0(n5597), .A1(n5016), .B0(n5598), .B1(n5020), .C0(n5599), 
        .C1(n5022), .Y(n6847) );
  MXI2X1 U8003 ( .A(\ImageBuffer[42][2] ), .B(n5013), .S0(n4896), .Y(n6849) );
  MXI2X1 U8004 ( .A(\ImageBuffer[41][2] ), .B(n5013), .S0(n4897), .Y(n6852) );
  OAI222XL U8005 ( .A0(n5615), .A1(n5016), .B0(n5616), .B1(n5020), .C0(n5617), 
        .C1(n5021), .Y(n6853) );
  MXI2X1 U8006 ( .A(\ImageBuffer[40][2] ), .B(n5013), .S0(n4898), .Y(n6855) );
  OAI222XL U8007 ( .A0(n5624), .A1(n5016), .B0(n5625), .B1(n5020), .C0(n5626), 
        .C1(n5024), .Y(n6856) );
  OAI21XL U8008 ( .A0(n6857), .A1(n5628), .B0(n6858), .Y(n8434) );
  MXI2X1 U8009 ( .A(\ImageBuffer[39][2] ), .B(n5013), .S0(n4900), .Y(n6858) );
  AOI211X1 U8010 ( .A0(n5082), .A1(n5631), .B0(n6859), .C0(n6785), .Y(n6857)
         );
  OAI222XL U8011 ( .A0(n5633), .A1(n5016), .B0(n5634), .B1(n5020), .C0(n5635), 
        .C1(n5023), .Y(n6859) );
  OAI21XL U8012 ( .A0(n6860), .A1(n5637), .B0(n6861), .Y(n8435) );
  MXI2X1 U8013 ( .A(\ImageBuffer[38][2] ), .B(n5013), .S0(n4901), .Y(n6861) );
  AOI211X1 U8014 ( .A0(n5082), .A1(n5640), .B0(n6862), .C0(n6785), .Y(n6860)
         );
  OAI222XL U8015 ( .A0(n5642), .A1(n5016), .B0(n5643), .B1(n5020), .C0(n5644), 
        .C1(n5022), .Y(n6862) );
  OAI21XL U8016 ( .A0(n6863), .A1(n5646), .B0(n6864), .Y(n8436) );
  MXI2X1 U8017 ( .A(\ImageBuffer[37][2] ), .B(n5013), .S0(n4902), .Y(n6864) );
  AOI211X1 U8018 ( .A0(n5082), .A1(n5649), .B0(n6865), .C0(n6785), .Y(n6863)
         );
  OAI222XL U8019 ( .A0(n5651), .A1(n5016), .B0(n5652), .B1(n5020), .C0(n5653), 
        .C1(n5023), .Y(n6865) );
  OAI21XL U8020 ( .A0(n6866), .A1(n5655), .B0(n6867), .Y(n8437) );
  MXI2X1 U8021 ( .A(\ImageBuffer[36][2] ), .B(n5013), .S0(n4903), .Y(n6867) );
  AOI211X1 U8022 ( .A0(n5082), .A1(n5658), .B0(n6868), .C0(n6785), .Y(n6866)
         );
  OAI222XL U8023 ( .A0(n5660), .A1(n5016), .B0(n5661), .B1(n5020), .C0(n5662), 
        .C1(n5022), .Y(n6868) );
  MXI2X1 U8024 ( .A(\ImageBuffer[35][2] ), .B(n5012), .S0(n4904), .Y(n6870) );
  OAI222XL U8025 ( .A0(n5669), .A1(n5015), .B0(n5670), .B1(n5020), .C0(n5671), 
        .C1(n5023), .Y(n6871) );
  MXI2X1 U8026 ( .A(\ImageBuffer[34][2] ), .B(n5012), .S0(n4905), .Y(n6873) );
  OAI222XL U8027 ( .A0(n5678), .A1(n5015), .B0(n5679), .B1(n5020), .C0(n5680), 
        .C1(n5023), .Y(n6874) );
  MXI2X1 U8028 ( .A(\ImageBuffer[33][2] ), .B(n5012), .S0(n4906), .Y(n6876) );
  OAI222XL U8029 ( .A0(n5687), .A1(n5015), .B0(n5688), .B1(n5020), .C0(n5689), 
        .C1(n5023), .Y(n6877) );
  MXI2X1 U8030 ( .A(\ImageBuffer[32][2] ), .B(n5012), .S0(n4907), .Y(n6879) );
  OAI222XL U8031 ( .A0(n5696), .A1(n5015), .B0(n5697), .B1(n5020), .C0(n5698), 
        .C1(n5023), .Y(n6880) );
  MXI2X1 U8032 ( .A(\ImageBuffer[31][2] ), .B(n5012), .S0(n4909), .Y(n6882) );
  OAI222XL U8033 ( .A0(n5705), .A1(n5015), .B0(n5706), .B1(n5020), .C0(n5707), 
        .C1(n5023), .Y(n6883) );
  MXI2X1 U8034 ( .A(\ImageBuffer[30][2] ), .B(n5012), .S0(n4910), .Y(n6885) );
  OAI222XL U8035 ( .A0(n5714), .A1(n5015), .B0(n5715), .B1(n5020), .C0(n5716), 
        .C1(n5023), .Y(n6886) );
  MXI2X1 U8036 ( .A(\ImageBuffer[29][2] ), .B(n5012), .S0(n4911), .Y(n6888) );
  MXI2X1 U8037 ( .A(\ImageBuffer[28][2] ), .B(n5012), .S0(n4912), .Y(n6891) );
  MXI2X1 U8038 ( .A(\ImageBuffer[27][2] ), .B(n5012), .S0(n4913), .Y(n6894) );
  OAI222XL U8039 ( .A0(n5741), .A1(n5015), .B0(n5742), .B1(n5019), .C0(n5743), 
        .C1(n5023), .Y(n6895) );
  OAI21XL U8040 ( .A0(n6896), .A1(n5745), .B0(n6897), .Y(n8447) );
  MXI2X1 U8041 ( .A(\ImageBuffer[26][2] ), .B(n5012), .S0(n4914), .Y(n6897) );
  AOI211X1 U8042 ( .A0(n5081), .A1(n5748), .B0(n6898), .C0(n6785), .Y(n6896)
         );
  OAI222XL U8043 ( .A0(n5750), .A1(n5015), .B0(n5751), .B1(n5020), .C0(n5752), 
        .C1(n5023), .Y(n6898) );
  MXI2X1 U8044 ( .A(\ImageBuffer[25][2] ), .B(n5012), .S0(n4915), .Y(n6900) );
  MXI2X1 U8045 ( .A(\ImageBuffer[24][2] ), .B(n5012), .S0(n4916), .Y(n6903) );
  OAI21XL U8046 ( .A0(n6905), .A1(n5772), .B0(n6906), .Y(n8450) );
  MXI2X1 U8047 ( .A(\ImageBuffer[23][2] ), .B(n5011), .S0(n4918), .Y(n6906) );
  AOI211X1 U8048 ( .A0(n5081), .A1(n5775), .B0(n6907), .C0(n6785), .Y(n6905)
         );
  OAI222XL U8049 ( .A0(n5777), .A1(n5016), .B0(n5778), .B1(n5018), .C0(n5779), 
        .C1(n5022), .Y(n6907) );
  OAI21XL U8050 ( .A0(n6908), .A1(n5781), .B0(n6909), .Y(n8451) );
  MXI2X1 U8051 ( .A(\ImageBuffer[22][2] ), .B(n5011), .S0(n4919), .Y(n6909) );
  AOI211X1 U8052 ( .A0(n5081), .A1(n5784), .B0(n6910), .C0(n6785), .Y(n6908)
         );
  OAI222XL U8053 ( .A0(n5786), .A1(n5015), .B0(n5787), .B1(n5018), .C0(n5788), 
        .C1(n5022), .Y(n6910) );
  OAI21XL U8054 ( .A0(n6911), .A1(n5790), .B0(n6912), .Y(n8452) );
  MXI2X1 U8055 ( .A(\ImageBuffer[21][2] ), .B(n5011), .S0(n4920), .Y(n6912) );
  AOI211X1 U8056 ( .A0(n5081), .A1(n5793), .B0(n6913), .C0(n6785), .Y(n6911)
         );
  OAI222XL U8057 ( .A0(n5795), .A1(n5016), .B0(n5796), .B1(n5018), .C0(n5797), 
        .C1(n5022), .Y(n6913) );
  OAI21XL U8058 ( .A0(n6914), .A1(n5799), .B0(n6915), .Y(n8453) );
  MXI2X1 U8059 ( .A(\ImageBuffer[20][2] ), .B(n5011), .S0(n4921), .Y(n6915) );
  AOI211X1 U8060 ( .A0(n5081), .A1(n5802), .B0(n6916), .C0(n6785), .Y(n6914)
         );
  OAI222XL U8061 ( .A0(n5804), .A1(n5016), .B0(n5805), .B1(n5018), .C0(n5806), 
        .C1(n5022), .Y(n6916) );
  MXI2X1 U8062 ( .A(\ImageBuffer[19][2] ), .B(n5011), .S0(n4922), .Y(n6918) );
  AOI211X1 U8063 ( .A0(n5081), .A1(n5811), .B0(n6919), .C0(n6785), .Y(n6917)
         );
  OAI222XL U8064 ( .A0(n5813), .A1(n5016), .B0(n5814), .B1(n5018), .C0(n5815), 
        .C1(n5022), .Y(n6919) );
  OAI21XL U8065 ( .A0(n6920), .A1(n5817), .B0(n6921), .Y(n8455) );
  MXI2X1 U8066 ( .A(\ImageBuffer[18][2] ), .B(n5011), .S0(n4923), .Y(n6921) );
  AOI211X1 U8067 ( .A0(n5081), .A1(n5820), .B0(n6922), .C0(n6785), .Y(n6920)
         );
  OAI222XL U8068 ( .A0(n5822), .A1(n5015), .B0(n5823), .B1(n5018), .C0(n5824), 
        .C1(n5022), .Y(n6922) );
  OAI21XL U8069 ( .A0(n6923), .A1(n5826), .B0(n6924), .Y(n8456) );
  MXI2X1 U8070 ( .A(\ImageBuffer[17][2] ), .B(n5011), .S0(n4924), .Y(n6924) );
  AOI211X1 U8071 ( .A0(n5081), .A1(n5829), .B0(n6925), .C0(n6785), .Y(n6923)
         );
  OAI222XL U8072 ( .A0(n5831), .A1(n5016), .B0(n5832), .B1(n5018), .C0(n5833), 
        .C1(n5022), .Y(n6925) );
  MXI2X1 U8073 ( .A(\ImageBuffer[16][2] ), .B(n5011), .S0(n4925), .Y(n6927) );
  OAI222XL U8074 ( .A0(n5840), .A1(n5015), .B0(n5841), .B1(n5018), .C0(n5842), 
        .C1(n5022), .Y(n6928) );
  OAI21XL U8075 ( .A0(n6929), .A1(n5844), .B0(n6930), .Y(n8458) );
  MXI2X1 U8076 ( .A(\ImageBuffer[15][2] ), .B(n5011), .S0(n4927), .Y(n6930) );
  AOI211X1 U8077 ( .A0(n5081), .A1(n5847), .B0(n6931), .C0(n6785), .Y(n6929)
         );
  OAI222XL U8078 ( .A0(n5849), .A1(n5017), .B0(n5850), .B1(n5018), .C0(n5851), 
        .C1(n5022), .Y(n6931) );
  OAI21XL U8079 ( .A0(n6932), .A1(n5853), .B0(n6933), .Y(n8459) );
  MXI2X1 U8080 ( .A(\ImageBuffer[14][2] ), .B(n5011), .S0(n4928), .Y(n6933) );
  AOI211X1 U8081 ( .A0(n5081), .A1(n5856), .B0(n6934), .C0(n6785), .Y(n6932)
         );
  OAI222XL U8082 ( .A0(n5858), .A1(n5015), .B0(n5859), .B1(n5018), .C0(n5860), 
        .C1(n5022), .Y(n6934) );
  OAI21XL U8083 ( .A0(n6935), .A1(n5862), .B0(n6936), .Y(n8460) );
  MXI2X1 U8084 ( .A(\ImageBuffer[13][2] ), .B(n5011), .S0(n4929), .Y(n6936) );
  AOI211X1 U8085 ( .A0(n5081), .A1(n5865), .B0(n6937), .C0(n6785), .Y(n6935)
         );
  OAI222XL U8086 ( .A0(n5867), .A1(n5016), .B0(n5868), .B1(n5018), .C0(n5869), 
        .C1(n5022), .Y(n6937) );
  MXI2X1 U8087 ( .A(\ImageBuffer[12][2] ), .B(n5011), .S0(n4930), .Y(n6939) );
  OAI222XL U8088 ( .A0(n5876), .A1(n5017), .B0(n5877), .B1(n5018), .C0(n5878), 
        .C1(n5022), .Y(n6940) );
  OAI21XL U8089 ( .A0(n6941), .A1(n5880), .B0(n6942), .Y(n8462) );
  MXI2X1 U8090 ( .A(\ImageBuffer[11][2] ), .B(n5011), .S0(n4931), .Y(n6942) );
  AOI211X1 U8091 ( .A0(n5081), .A1(n5883), .B0(n6943), .C0(n6785), .Y(n6941)
         );
  OAI222XL U8092 ( .A0(n5885), .A1(n6786), .B0(n5886), .B1(n5019), .C0(n5887), 
        .C1(n5021), .Y(n6943) );
  OAI21XL U8093 ( .A0(n6944), .A1(n5889), .B0(n6945), .Y(n8463) );
  MXI2X1 U8094 ( .A(\ImageBuffer[10][2] ), .B(n5014), .S0(n4932), .Y(n6945) );
  AOI211X1 U8095 ( .A0(n5081), .A1(n5892), .B0(n6946), .C0(n6785), .Y(n6944)
         );
  OAI222XL U8096 ( .A0(n5894), .A1(n6786), .B0(n5895), .B1(n5019), .C0(n5896), 
        .C1(n5021), .Y(n6946) );
  OAI21XL U8097 ( .A0(n6947), .A1(n5898), .B0(n6948), .Y(n8464) );
  MXI2X1 U8098 ( .A(\ImageBuffer[9][2] ), .B(n5013), .S0(n4933), .Y(n6948) );
  AOI211X1 U8099 ( .A0(n5081), .A1(n5901), .B0(n6949), .C0(n6785), .Y(n6947)
         );
  OAI222XL U8100 ( .A0(n5903), .A1(n5016), .B0(n5904), .B1(n5019), .C0(n5905), 
        .C1(n5021), .Y(n6949) );
  OAI21XL U8101 ( .A0(n6950), .A1(n5907), .B0(n6951), .Y(n8465) );
  MXI2X1 U8102 ( .A(\ImageBuffer[8][2] ), .B(n5012), .S0(n4934), .Y(n6951) );
  AOI211X1 U8103 ( .A0(n5081), .A1(n5910), .B0(n6952), .C0(n6785), .Y(n6950)
         );
  OAI222XL U8104 ( .A0(n5912), .A1(n5015), .B0(n5913), .B1(n5019), .C0(n5914), 
        .C1(n5021), .Y(n6952) );
  OAI21XL U8105 ( .A0(n6953), .A1(n5916), .B0(n6954), .Y(n8466) );
  MXI2X1 U8106 ( .A(\ImageBuffer[7][2] ), .B(n5011), .S0(n4935), .Y(n6954) );
  AOI211X1 U8107 ( .A0(n5081), .A1(n5919), .B0(n6955), .C0(n6785), .Y(n6953)
         );
  OAI222XL U8108 ( .A0(n5921), .A1(n5017), .B0(n5922), .B1(n5019), .C0(n5923), 
        .C1(n5021), .Y(n6955) );
  OAI21XL U8109 ( .A0(n6956), .A1(n5925), .B0(n6957), .Y(n8467) );
  MXI2X1 U8110 ( .A(\ImageBuffer[6][2] ), .B(n5014), .S0(n4936), .Y(n6957) );
  AOI211X1 U8111 ( .A0(n5081), .A1(n5928), .B0(n6958), .C0(n6785), .Y(n6956)
         );
  OAI222XL U8112 ( .A0(n5930), .A1(n5015), .B0(n5931), .B1(n5019), .C0(n5932), 
        .C1(n5021), .Y(n6958) );
  OAI21XL U8113 ( .A0(n6959), .A1(n5934), .B0(n6960), .Y(n8468) );
  MXI2X1 U8114 ( .A(\ImageBuffer[5][2] ), .B(n5013), .S0(n4937), .Y(n6960) );
  AOI211X1 U8115 ( .A0(n5081), .A1(n5937), .B0(n6961), .C0(n6785), .Y(n6959)
         );
  OAI222XL U8116 ( .A0(n5939), .A1(n5016), .B0(n5940), .B1(n5019), .C0(n5941), 
        .C1(n5021), .Y(n6961) );
  OAI21XL U8117 ( .A0(n6962), .A1(n5943), .B0(n6963), .Y(n8469) );
  MXI2X1 U8118 ( .A(\ImageBuffer[4][2] ), .B(n5014), .S0(n4938), .Y(n6963) );
  AOI211X1 U8119 ( .A0(n5081), .A1(n5946), .B0(n6964), .C0(n6785), .Y(n6962)
         );
  OAI222XL U8120 ( .A0(n5948), .A1(n5015), .B0(n5949), .B1(n5019), .C0(n5950), 
        .C1(n5021), .Y(n6964) );
  OAI21XL U8121 ( .A0(n6965), .A1(n5952), .B0(n6966), .Y(n8470) );
  MXI2X1 U8122 ( .A(\ImageBuffer[3][2] ), .B(n5013), .S0(n4939), .Y(n6966) );
  AOI211X1 U8123 ( .A0(n5081), .A1(n5955), .B0(n6967), .C0(n6785), .Y(n6965)
         );
  OAI222XL U8124 ( .A0(n5957), .A1(n5017), .B0(n5958), .B1(n5019), .C0(n5959), 
        .C1(n5021), .Y(n6967) );
  MXI2X1 U8125 ( .A(\ImageBuffer[2][2] ), .B(n5014), .S0(n4940), .Y(n6969) );
  OAI21XL U8126 ( .A0(n6971), .A1(n5970), .B0(n6972), .Y(n8472) );
  MXI2X1 U8127 ( .A(\ImageBuffer[1][2] ), .B(n5013), .S0(n4941), .Y(n6972) );
  AOI211X1 U8128 ( .A0(n5081), .A1(n5973), .B0(n6973), .C0(n6785), .Y(n6971)
         );
  OAI222XL U8129 ( .A0(n5975), .A1(n6786), .B0(n5976), .B1(n5019), .C0(n5977), 
        .C1(n5021), .Y(n6973) );
  MXI2X1 U8130 ( .A(\ImageBuffer[0][2] ), .B(n5014), .S0(n4942), .Y(n6975) );
  NOR2BX1 U8131 ( .AN(IROM_Q[2]), .B(n4945), .Y(n6783) );
  AOI211X1 U8132 ( .A0(n5082), .A1(n5983), .B0(n6976), .C0(n6785), .Y(n6974)
         );
  OAI222XL U8133 ( .A0(n5989), .A1(n5015), .B0(n5990), .B1(n5019), .C0(n5991), 
        .C1(n5021), .Y(n6976) );
  CLKINVX1 U8134 ( .A(n4872), .Y(n6786) );
  OAI21XL U8135 ( .A0(n6978), .A1(n5408), .B0(n6979), .Y(n8474) );
  AOI211X1 U8136 ( .A0(n5077), .A1(n5412), .B0(n6981), .C0(n6982), .Y(n6978)
         );
  OAI222XL U8137 ( .A0(n5415), .A1(n5030), .B0(n5416), .B1(n5033), .C0(n5418), 
        .C1(n5036), .Y(n6981) );
  OAI21XL U8138 ( .A0(n6986), .A1(n5421), .B0(n6987), .Y(n8475) );
  OAI222XL U8139 ( .A0(n5426), .A1(n5030), .B0(n5427), .B1(n5032), .C0(n5428), 
        .C1(n5036), .Y(n6988) );
  OAI21XL U8140 ( .A0(n6989), .A1(n5430), .B0(n6990), .Y(n8476) );
  OAI222XL U8141 ( .A0(n5435), .A1(n5030), .B0(n5436), .B1(n5031), .C0(n5437), 
        .C1(n5036), .Y(n6991) );
  OAI21XL U8142 ( .A0(n6992), .A1(n5439), .B0(n6993), .Y(n8477) );
  OAI222XL U8143 ( .A0(n5444), .A1(n5030), .B0(n5445), .B1(n5034), .C0(n5446), 
        .C1(n5036), .Y(n6994) );
  OAI21XL U8144 ( .A0(n6995), .A1(n5448), .B0(n6996), .Y(n8478) );
  OAI222XL U8145 ( .A0(n5453), .A1(n5028), .B0(n5454), .B1(n5034), .C0(n5455), 
        .C1(n5036), .Y(n6997) );
  OAI21XL U8146 ( .A0(n6998), .A1(n5457), .B0(n6999), .Y(n8479) );
  MXI2X1 U8147 ( .A(\ImageBuffer[58][1] ), .B(n5027), .S0(n4878), .Y(n6999) );
  OAI222XL U8148 ( .A0(n5462), .A1(n5028), .B0(n5463), .B1(n5034), .C0(n5464), 
        .C1(n5037), .Y(n7000) );
  OAI21XL U8149 ( .A0(n7001), .A1(n5466), .B0(n7002), .Y(n8480) );
  OAI222XL U8150 ( .A0(n5471), .A1(n5028), .B0(n5472), .B1(n5034), .C0(n5473), 
        .C1(n5037), .Y(n7003) );
  OAI21XL U8151 ( .A0(n7004), .A1(n5475), .B0(n7005), .Y(n8481) );
  MXI2X1 U8152 ( .A(\ImageBuffer[56][1] ), .B(n5027), .S0(n4880), .Y(n7005) );
  AOI211X1 U8153 ( .A0(n5076), .A1(n5478), .B0(n7006), .C0(n6982), .Y(n7004)
         );
  OAI222XL U8154 ( .A0(n5480), .A1(n6983), .B0(n5481), .B1(n5034), .C0(n5482), 
        .C1(n5037), .Y(n7006) );
  OAI21XL U8155 ( .A0(n7007), .A1(n5484), .B0(n7008), .Y(n8482) );
  AOI211X1 U8156 ( .A0(n5076), .A1(n5487), .B0(n7009), .C0(n6982), .Y(n7007)
         );
  OAI222XL U8157 ( .A0(n5489), .A1(n5028), .B0(n5490), .B1(n5034), .C0(n5491), 
        .C1(n5037), .Y(n7009) );
  OAI21XL U8158 ( .A0(n7010), .A1(n5493), .B0(n7011), .Y(n8483) );
  AOI211X1 U8159 ( .A0(n5076), .A1(n5496), .B0(n7012), .C0(n6982), .Y(n7010)
         );
  OAI21XL U8160 ( .A0(n7013), .A1(n5502), .B0(n7014), .Y(n8484) );
  AOI211X1 U8161 ( .A0(n5076), .A1(n5505), .B0(n7015), .C0(n6982), .Y(n7013)
         );
  OAI222XL U8162 ( .A0(n5507), .A1(n5028), .B0(n5508), .B1(n5034), .C0(n5509), 
        .C1(n5037), .Y(n7015) );
  OAI21XL U8163 ( .A0(n7016), .A1(n5511), .B0(n7017), .Y(n8485) );
  OAI222XL U8164 ( .A0(n5516), .A1(n5028), .B0(n5517), .B1(n5034), .C0(n5518), 
        .C1(n5037), .Y(n7018) );
  OAI21XL U8165 ( .A0(n7019), .A1(n5520), .B0(n7020), .Y(n8486) );
  AOI211X1 U8166 ( .A0(n5076), .A1(n5523), .B0(n7021), .C0(n6982), .Y(n7019)
         );
  OAI222XL U8167 ( .A0(n5525), .A1(n5030), .B0(n5526), .B1(n5034), .C0(n5527), 
        .C1(n5035), .Y(n7021) );
  OAI21XL U8168 ( .A0(n7022), .A1(n5529), .B0(n7023), .Y(n8487) );
  MXI2X1 U8169 ( .A(\ImageBuffer[50][1] ), .B(n5027), .S0(n4887), .Y(n7023) );
  AOI211X1 U8170 ( .A0(n5076), .A1(n5532), .B0(n7024), .C0(n6982), .Y(n7022)
         );
  OAI222XL U8171 ( .A0(n5534), .A1(n6983), .B0(n5535), .B1(n5034), .C0(n5536), 
        .C1(n5035), .Y(n7024) );
  OAI21XL U8172 ( .A0(n7025), .A1(n5538), .B0(n7026), .Y(n8488) );
  OAI222XL U8173 ( .A0(n5543), .A1(n5028), .B0(n5544), .B1(n5034), .C0(n5545), 
        .C1(n5036), .Y(n7027) );
  OAI21XL U8174 ( .A0(n7028), .A1(n5547), .B0(n7029), .Y(n8489) );
  AOI211X1 U8175 ( .A0(n5076), .A1(n5550), .B0(n7030), .C0(n6982), .Y(n7028)
         );
  OAI222XL U8176 ( .A0(n5552), .A1(n6983), .B0(n5553), .B1(n5034), .C0(n5554), 
        .C1(n5035), .Y(n7030) );
  OAI21XL U8177 ( .A0(n7031), .A1(n5556), .B0(n7032), .Y(n8490) );
  AOI211X1 U8178 ( .A0(n5076), .A1(n5559), .B0(n7033), .C0(n6982), .Y(n7031)
         );
  OAI222XL U8179 ( .A0(n5561), .A1(n5029), .B0(n5562), .B1(n5033), .C0(n5563), 
        .C1(n5037), .Y(n7033) );
  OAI21XL U8180 ( .A0(n7034), .A1(n5565), .B0(n7035), .Y(n8491) );
  MXI2X1 U8181 ( .A(\ImageBuffer[46][1] ), .B(n5026), .S0(n4892), .Y(n7035) );
  AOI211X1 U8182 ( .A0(n5076), .A1(n5568), .B0(n7036), .C0(n6982), .Y(n7034)
         );
  OAI222XL U8183 ( .A0(n5570), .A1(n5029), .B0(n5571), .B1(n5033), .C0(n5572), 
        .C1(n5037), .Y(n7036) );
  OAI21XL U8184 ( .A0(n7037), .A1(n5574), .B0(n7038), .Y(n8492) );
  AOI211X1 U8185 ( .A0(n5076), .A1(n5577), .B0(n7039), .C0(n6982), .Y(n7037)
         );
  OAI222XL U8186 ( .A0(n5579), .A1(n5028), .B0(n5580), .B1(n5033), .C0(n5581), 
        .C1(n5037), .Y(n7039) );
  OAI21XL U8187 ( .A0(n7040), .A1(n5583), .B0(n7041), .Y(n8493) );
  MXI2X1 U8188 ( .A(\ImageBuffer[44][1] ), .B(n5026), .S0(n4894), .Y(n7041) );
  AOI211X1 U8189 ( .A0(n5076), .A1(n5586), .B0(n7042), .C0(n6982), .Y(n7040)
         );
  OAI222XL U8190 ( .A0(n5588), .A1(n5029), .B0(n5589), .B1(n5033), .C0(n5590), 
        .C1(n5037), .Y(n7042) );
  OAI21XL U8191 ( .A0(n7043), .A1(n5592), .B0(n7044), .Y(n8494) );
  AOI211X1 U8192 ( .A0(n5076), .A1(n5595), .B0(n7045), .C0(n6982), .Y(n7043)
         );
  OAI222XL U8193 ( .A0(n5597), .A1(n5028), .B0(n5598), .B1(n5033), .C0(n5599), 
        .C1(n5037), .Y(n7045) );
  OAI21XL U8194 ( .A0(n7046), .A1(n5601), .B0(n7047), .Y(n8495) );
  AOI211X1 U8195 ( .A0(n5076), .A1(n5604), .B0(n7048), .C0(n6982), .Y(n7046)
         );
  OAI222XL U8196 ( .A0(n5606), .A1(n5029), .B0(n5607), .B1(n5033), .C0(n5608), 
        .C1(n5037), .Y(n7048) );
  OAI21XL U8197 ( .A0(n7049), .A1(n5610), .B0(n7050), .Y(n8496) );
  AOI211X1 U8198 ( .A0(n5076), .A1(n5613), .B0(n7051), .C0(n6982), .Y(n7049)
         );
  OAI222XL U8199 ( .A0(n5615), .A1(n5028), .B0(n5616), .B1(n5033), .C0(n5617), 
        .C1(n5037), .Y(n7051) );
  OAI21XL U8200 ( .A0(n7052), .A1(n5619), .B0(n7053), .Y(n8497) );
  AOI211X1 U8201 ( .A0(n5076), .A1(n5622), .B0(n7054), .C0(n6982), .Y(n7052)
         );
  OAI222XL U8202 ( .A0(n5624), .A1(n5029), .B0(n5625), .B1(n5033), .C0(n5626), 
        .C1(n5037), .Y(n7054) );
  OAI21XL U8203 ( .A0(n7055), .A1(n5628), .B0(n7056), .Y(n8498) );
  AOI211X1 U8204 ( .A0(n5076), .A1(n5631), .B0(n7057), .C0(n6982), .Y(n7055)
         );
  OAI222XL U8205 ( .A0(n5633), .A1(n5029), .B0(n5634), .B1(n5033), .C0(n5635), 
        .C1(n5037), .Y(n7057) );
  OAI21XL U8206 ( .A0(n7058), .A1(n5637), .B0(n7059), .Y(n8499) );
  AOI211X1 U8207 ( .A0(n5076), .A1(n5640), .B0(n7060), .C0(n6982), .Y(n7058)
         );
  OAI222XL U8208 ( .A0(n5642), .A1(n5028), .B0(n5643), .B1(n5033), .C0(n5644), 
        .C1(n5037), .Y(n7060) );
  OAI21XL U8209 ( .A0(n7061), .A1(n5646), .B0(n7062), .Y(n8500) );
  AOI211X1 U8210 ( .A0(n5076), .A1(n5649), .B0(n7063), .C0(n6982), .Y(n7061)
         );
  OAI222XL U8211 ( .A0(n5651), .A1(n5028), .B0(n5652), .B1(n5033), .C0(n5653), 
        .C1(n5037), .Y(n7063) );
  OAI21XL U8212 ( .A0(n7064), .A1(n5655), .B0(n7065), .Y(n8501) );
  AOI211X1 U8213 ( .A0(n5076), .A1(n5658), .B0(n7066), .C0(n6982), .Y(n7064)
         );
  OAI222XL U8214 ( .A0(n5660), .A1(n5029), .B0(n5661), .B1(n5033), .C0(n5662), 
        .C1(n5037), .Y(n7066) );
  OAI21XL U8215 ( .A0(n7067), .A1(n5664), .B0(n7068), .Y(n8502) );
  AOI211X1 U8216 ( .A0(n5076), .A1(n5667), .B0(n7069), .C0(n6982), .Y(n7067)
         );
  OAI222XL U8217 ( .A0(n5669), .A1(n5028), .B0(n5670), .B1(n5034), .C0(n5671), 
        .C1(n5035), .Y(n7069) );
  OAI21XL U8218 ( .A0(n7070), .A1(n5673), .B0(n7071), .Y(n8503) );
  AOI211X1 U8219 ( .A0(n5076), .A1(n5676), .B0(n7072), .C0(n6982), .Y(n7070)
         );
  OAI222XL U8220 ( .A0(n5678), .A1(n5029), .B0(n5679), .B1(n5034), .C0(n5680), 
        .C1(n5035), .Y(n7072) );
  OAI21XL U8221 ( .A0(n7073), .A1(n5682), .B0(n7074), .Y(n8504) );
  AOI211X1 U8222 ( .A0(n5076), .A1(n5685), .B0(n7075), .C0(n6982), .Y(n7073)
         );
  OAI222XL U8223 ( .A0(n5687), .A1(n5028), .B0(n5688), .B1(n5031), .C0(n5689), 
        .C1(n5036), .Y(n7075) );
  OAI21XL U8224 ( .A0(n7076), .A1(n5691), .B0(n7077), .Y(n8505) );
  AOI211X1 U8225 ( .A0(n5076), .A1(n5694), .B0(n7078), .C0(n6982), .Y(n7076)
         );
  OAI222XL U8226 ( .A0(n5696), .A1(n5030), .B0(n5697), .B1(n5034), .C0(n5698), 
        .C1(n5035), .Y(n7078) );
  OAI21XL U8227 ( .A0(n7079), .A1(n5700), .B0(n7080), .Y(n8506) );
  AOI211X1 U8228 ( .A0(n5076), .A1(n5703), .B0(n7081), .C0(n6982), .Y(n7079)
         );
  OAI222XL U8229 ( .A0(n5705), .A1(n5029), .B0(n5706), .B1(n5031), .C0(n5707), 
        .C1(n5035), .Y(n7081) );
  OAI21XL U8230 ( .A0(n7082), .A1(n5709), .B0(n7083), .Y(n8507) );
  AOI211X1 U8231 ( .A0(n5076), .A1(n5712), .B0(n7084), .C0(n6982), .Y(n7082)
         );
  OAI222XL U8232 ( .A0(n5714), .A1(n5030), .B0(n5715), .B1(n5031), .C0(n5716), 
        .C1(n5036), .Y(n7084) );
  OAI21XL U8233 ( .A0(n7085), .A1(n5718), .B0(n7086), .Y(n8508) );
  AOI211X1 U8234 ( .A0(n5076), .A1(n5721), .B0(n7087), .C0(n6982), .Y(n7085)
         );
  OAI222XL U8235 ( .A0(n5723), .A1(n5030), .B0(n5724), .B1(n5034), .C0(n5725), 
        .C1(n5035), .Y(n7087) );
  OAI21XL U8236 ( .A0(n7088), .A1(n5727), .B0(n7089), .Y(n8509) );
  AOI211X1 U8237 ( .A0(n5076), .A1(n5730), .B0(n7090), .C0(n6982), .Y(n7088)
         );
  OAI222XL U8238 ( .A0(n5732), .A1(n5030), .B0(n5733), .B1(n5031), .C0(n5734), 
        .C1(n5035), .Y(n7090) );
  OAI21XL U8239 ( .A0(n7091), .A1(n5736), .B0(n7092), .Y(n8510) );
  AOI211X1 U8240 ( .A0(n5075), .A1(n5739), .B0(n7093), .C0(n6982), .Y(n7091)
         );
  OAI222XL U8241 ( .A0(n5741), .A1(n5028), .B0(n5742), .B1(n5034), .C0(n5743), 
        .C1(n5035), .Y(n7093) );
  OAI21XL U8242 ( .A0(n7094), .A1(n5745), .B0(n7095), .Y(n8511) );
  AOI211X1 U8243 ( .A0(n5075), .A1(n5748), .B0(n7096), .C0(n6982), .Y(n7094)
         );
  OAI21XL U8244 ( .A0(n7097), .A1(n5754), .B0(n7098), .Y(n8512) );
  AOI211X1 U8245 ( .A0(n5075), .A1(n5757), .B0(n7099), .C0(n6982), .Y(n7097)
         );
  OAI222XL U8246 ( .A0(n5759), .A1(n6983), .B0(n5760), .B1(n5031), .C0(n5761), 
        .C1(n6985), .Y(n7099) );
  OAI21XL U8247 ( .A0(n7100), .A1(n5763), .B0(n7101), .Y(n8513) );
  AOI211X1 U8248 ( .A0(n5075), .A1(n5766), .B0(n7102), .C0(n6982), .Y(n7100)
         );
  OAI222XL U8249 ( .A0(n5768), .A1(n5028), .B0(n5769), .B1(n5031), .C0(n5770), 
        .C1(n5035), .Y(n7102) );
  OAI21XL U8250 ( .A0(n7103), .A1(n5772), .B0(n7104), .Y(n8514) );
  AOI211X1 U8251 ( .A0(n5075), .A1(n5775), .B0(n7105), .C0(n6982), .Y(n7103)
         );
  OAI222XL U8252 ( .A0(n5777), .A1(n5030), .B0(n5778), .B1(n5032), .C0(n5779), 
        .C1(n5036), .Y(n7105) );
  OAI21XL U8253 ( .A0(n7106), .A1(n5781), .B0(n7107), .Y(n8515) );
  AOI211X1 U8254 ( .A0(n5075), .A1(n5784), .B0(n7108), .C0(n6982), .Y(n7106)
         );
  OAI222XL U8255 ( .A0(n5786), .A1(n5030), .B0(n5787), .B1(n5032), .C0(n5788), 
        .C1(n5036), .Y(n7108) );
  OAI21XL U8256 ( .A0(n7109), .A1(n5790), .B0(n7110), .Y(n8516) );
  AOI211X1 U8257 ( .A0(n5075), .A1(n5793), .B0(n7111), .C0(n6982), .Y(n7109)
         );
  OAI222XL U8258 ( .A0(n5795), .A1(n5030), .B0(n5796), .B1(n5032), .C0(n5797), 
        .C1(n5036), .Y(n7111) );
  OAI21XL U8259 ( .A0(n7112), .A1(n5799), .B0(n7113), .Y(n8517) );
  AOI211X1 U8260 ( .A0(n5075), .A1(n5802), .B0(n7114), .C0(n6982), .Y(n7112)
         );
  OAI222XL U8261 ( .A0(n5804), .A1(n5030), .B0(n5805), .B1(n5032), .C0(n5806), 
        .C1(n5036), .Y(n7114) );
  OAI21XL U8262 ( .A0(n7115), .A1(n5808), .B0(n7116), .Y(n8518) );
  MXI2X1 U8263 ( .A(\ImageBuffer[19][1] ), .B(n5025), .S0(n4922), .Y(n7116) );
  AOI211X1 U8264 ( .A0(n5075), .A1(n5811), .B0(n7117), .C0(n6982), .Y(n7115)
         );
  OAI222XL U8265 ( .A0(n5813), .A1(n5030), .B0(n5814), .B1(n5032), .C0(n5815), 
        .C1(n5036), .Y(n7117) );
  OAI21XL U8266 ( .A0(n7118), .A1(n5817), .B0(n7119), .Y(n8519) );
  AOI211X1 U8267 ( .A0(n5075), .A1(n5820), .B0(n7120), .C0(n6982), .Y(n7118)
         );
  OAI222XL U8268 ( .A0(n5822), .A1(n5030), .B0(n5823), .B1(n5032), .C0(n5824), 
        .C1(n5036), .Y(n7120) );
  OAI21XL U8269 ( .A0(n7121), .A1(n5826), .B0(n7122), .Y(n8520) );
  AOI211X1 U8270 ( .A0(n5075), .A1(n5829), .B0(n7123), .C0(n6982), .Y(n7121)
         );
  OAI222XL U8271 ( .A0(n5831), .A1(n5030), .B0(n5832), .B1(n5032), .C0(n5833), 
        .C1(n5036), .Y(n7123) );
  OAI21XL U8272 ( .A0(n7124), .A1(n5835), .B0(n7125), .Y(n8521) );
  MXI2X1 U8273 ( .A(\ImageBuffer[16][1] ), .B(n5025), .S0(n4925), .Y(n7125) );
  AOI211X1 U8274 ( .A0(n5075), .A1(n5838), .B0(n7126), .C0(n6982), .Y(n7124)
         );
  OAI222XL U8275 ( .A0(n5840), .A1(n5030), .B0(n5841), .B1(n5032), .C0(n5842), 
        .C1(n5036), .Y(n7126) );
  OAI21XL U8276 ( .A0(n7127), .A1(n5844), .B0(n7128), .Y(n8522) );
  AOI211X1 U8277 ( .A0(n5075), .A1(n5847), .B0(n7129), .C0(n6982), .Y(n7127)
         );
  OAI222XL U8278 ( .A0(n5849), .A1(n5030), .B0(n5850), .B1(n5032), .C0(n5851), 
        .C1(n5036), .Y(n7129) );
  OAI21XL U8279 ( .A0(n7130), .A1(n5853), .B0(n7131), .Y(n8523) );
  AOI211X1 U8280 ( .A0(n5075), .A1(n5856), .B0(n7132), .C0(n6982), .Y(n7130)
         );
  OAI222XL U8281 ( .A0(n5858), .A1(n5030), .B0(n5859), .B1(n5032), .C0(n5860), 
        .C1(n5036), .Y(n7132) );
  OAI21XL U8282 ( .A0(n7133), .A1(n5862), .B0(n7134), .Y(n8524) );
  AOI211X1 U8283 ( .A0(n5075), .A1(n5865), .B0(n7135), .C0(n6982), .Y(n7133)
         );
  OAI222XL U8284 ( .A0(n5867), .A1(n5030), .B0(n5868), .B1(n5032), .C0(n5869), 
        .C1(n5036), .Y(n7135) );
  OAI21XL U8285 ( .A0(n7136), .A1(n5871), .B0(n7137), .Y(n8525) );
  AOI211X1 U8286 ( .A0(n5075), .A1(n5874), .B0(n7138), .C0(n6982), .Y(n7136)
         );
  OAI222XL U8287 ( .A0(n5876), .A1(n5030), .B0(n5877), .B1(n5032), .C0(n5878), 
        .C1(n5036), .Y(n7138) );
  OAI21XL U8288 ( .A0(n7139), .A1(n5880), .B0(n7140), .Y(n8526) );
  AOI211X1 U8289 ( .A0(n5075), .A1(n5883), .B0(n7141), .C0(n6982), .Y(n7139)
         );
  OAI222XL U8290 ( .A0(n5885), .A1(n5029), .B0(n5886), .B1(n5031), .C0(n5887), 
        .C1(n5035), .Y(n7141) );
  OAI21XL U8291 ( .A0(n7142), .A1(n5889), .B0(n7143), .Y(n8527) );
  AOI211X1 U8292 ( .A0(n5075), .A1(n5892), .B0(n7144), .C0(n6982), .Y(n7142)
         );
  OAI222XL U8293 ( .A0(n5894), .A1(n5029), .B0(n5895), .B1(n5031), .C0(n5896), 
        .C1(n5037), .Y(n7144) );
  OAI21XL U8294 ( .A0(n7145), .A1(n5898), .B0(n7146), .Y(n8528) );
  AOI211X1 U8295 ( .A0(n5075), .A1(n5901), .B0(n7147), .C0(n6982), .Y(n7145)
         );
  OAI222XL U8296 ( .A0(n5903), .A1(n5029), .B0(n5904), .B1(n5031), .C0(n5905), 
        .C1(n5155), .Y(n7147) );
  OAI21XL U8297 ( .A0(n7148), .A1(n5907), .B0(n7149), .Y(n8529) );
  MXI2X1 U8298 ( .A(\ImageBuffer[8][1] ), .B(n5027), .S0(n4934), .Y(n7149) );
  AOI211X1 U8299 ( .A0(n5075), .A1(n5910), .B0(n7150), .C0(n6982), .Y(n7148)
         );
  OAI222XL U8300 ( .A0(n5912), .A1(n5029), .B0(n5913), .B1(n5031), .C0(n5914), 
        .C1(n5037), .Y(n7150) );
  OAI21XL U8301 ( .A0(n7151), .A1(n5916), .B0(n7152), .Y(n8530) );
  AOI211X1 U8302 ( .A0(n5075), .A1(n5919), .B0(n7153), .C0(n6982), .Y(n7151)
         );
  OAI222XL U8303 ( .A0(n5921), .A1(n5029), .B0(n5922), .B1(n5031), .C0(n5923), 
        .C1(n5037), .Y(n7153) );
  OAI21XL U8304 ( .A0(n7154), .A1(n5925), .B0(n7155), .Y(n8531) );
  AOI211X1 U8305 ( .A0(n5075), .A1(n5928), .B0(n7156), .C0(n6982), .Y(n7154)
         );
  OAI222XL U8306 ( .A0(n5930), .A1(n5029), .B0(n5931), .B1(n5031), .C0(n5932), 
        .C1(n5035), .Y(n7156) );
  OAI21XL U8307 ( .A0(n7157), .A1(n5934), .B0(n7158), .Y(n8532) );
  AOI211X1 U8308 ( .A0(n5075), .A1(n5937), .B0(n7159), .C0(n6982), .Y(n7157)
         );
  OAI222XL U8309 ( .A0(n5939), .A1(n5029), .B0(n5940), .B1(n5031), .C0(n5941), 
        .C1(n5036), .Y(n7159) );
  OAI21XL U8310 ( .A0(n7160), .A1(n5943), .B0(n7161), .Y(n8533) );
  AOI211X1 U8311 ( .A0(n5075), .A1(n5946), .B0(n7162), .C0(n6982), .Y(n7160)
         );
  OAI222XL U8312 ( .A0(n5948), .A1(n5029), .B0(n5949), .B1(n5031), .C0(n5950), 
        .C1(n5035), .Y(n7162) );
  OAI21XL U8313 ( .A0(n7163), .A1(n5952), .B0(n7164), .Y(n8534) );
  AOI211X1 U8314 ( .A0(n5075), .A1(n5955), .B0(n7165), .C0(n6982), .Y(n7163)
         );
  OAI222XL U8315 ( .A0(n5957), .A1(n5029), .B0(n5958), .B1(n5031), .C0(n5959), 
        .C1(n5035), .Y(n7165) );
  OAI21XL U8316 ( .A0(n7166), .A1(n5961), .B0(n7167), .Y(n8535) );
  AOI211X1 U8317 ( .A0(n5075), .A1(n5964), .B0(n7168), .C0(n6982), .Y(n7166)
         );
  OAI21XL U8318 ( .A0(n7169), .A1(n5970), .B0(n7170), .Y(n8536) );
  AOI211X1 U8319 ( .A0(n5075), .A1(n5973), .B0(n7171), .C0(n6982), .Y(n7169)
         );
  OAI222XL U8320 ( .A0(n5975), .A1(n5029), .B0(n5976), .B1(n5031), .C0(n5977), 
        .C1(n5035), .Y(n7171) );
  OAI21XL U8321 ( .A0(n7172), .A1(n5979), .B0(n7173), .Y(n8537) );
  MXI2X1 U8322 ( .A(\ImageBuffer[0][1] ), .B(n5026), .S0(n4942), .Y(n7173) );
  NOR2BX1 U8323 ( .AN(IROM_Q[1]), .B(n4945), .Y(n6980) );
  AOI211X1 U8324 ( .A0(n5076), .A1(n5983), .B0(n7174), .C0(n6982), .Y(n7172)
         );
  OAI222XL U8325 ( .A0(n5989), .A1(n5029), .B0(n5990), .B1(n5031), .C0(n5991), 
        .C1(n5035), .Y(n7174) );
  CLKINVX1 U8326 ( .A(n4873), .Y(n6983) );
  OAI21XL U8327 ( .A0(n7176), .A1(n5408), .B0(n7177), .Y(n8538) );
  MXI2X1 U8328 ( .A(\ImageBuffer[63][0] ), .B(n5040), .S0(n5411), .Y(n7177) );
  OAI32X1 U8329 ( .A0(n7184), .A1(n5056), .A2(n7185), .B0(n3352), .B1(n7198), 
        .Y(n7199) );
  CLKINVX1 U8330 ( .A(n7191), .Y(n7185) );
  NAND2X1 U8331 ( .A(n7203), .B(n7204), .Y(n7198) );
  OAI21XL U8332 ( .A0(n7205), .A1(n5421), .B0(n7206), .Y(n8539) );
  MXI2X1 U8333 ( .A(\ImageBuffer[62][0] ), .B(n5040), .S0(n4874), .Y(n7206) );
  AOI211X1 U8334 ( .A0(n7210), .A1(n7183), .B0(n7211), .C0(n7212), .Y(n7209)
         );
  CLKINVX1 U8335 ( .A(n7215), .Y(n7212) );
  CLKINVX1 U8336 ( .A(n7232), .Y(n7230) );
  CLKINVX1 U8337 ( .A(n7229), .Y(n7226) );
  NAND2X1 U8338 ( .A(n7235), .B(n7204), .Y(n7232) );
  AOI211X1 U8339 ( .A0(n7240), .A1(n7183), .B0(n7241), .C0(n7242), .Y(n7239)
         );
  CLKINVX1 U8340 ( .A(n7245), .Y(n7242) );
  OAI21XL U8341 ( .A0(n7251), .A1(n5448), .B0(n7252), .Y(n8542) );
  MXI2X1 U8342 ( .A(\ImageBuffer[59][0] ), .B(n5039), .S0(n4877), .Y(n7252) );
  CLKINVX1 U8343 ( .A(n7260), .Y(n7257) );
  MXI2X1 U8344 ( .A(\ImageBuffer[58][0] ), .B(n5039), .S0(n4878), .Y(n7265) );
  CLKINVX1 U8345 ( .A(n7275), .Y(n7273) );
  CLKINVX1 U8346 ( .A(n7272), .Y(n7269) );
  NAND2X1 U8347 ( .A(n7277), .B(n7204), .Y(n7275) );
  MXI2X1 U8348 ( .A(\ImageBuffer[57][0] ), .B(n5039), .S0(n4879), .Y(n7279) );
  CLKINVX1 U8349 ( .A(n7287), .Y(n7284) );
  OAI21XL U8350 ( .A0(n7291), .A1(n5475), .B0(n7292), .Y(n8545) );
  MXI2X1 U8351 ( .A(\ImageBuffer[56][0] ), .B(n5039), .S0(n4880), .Y(n7292) );
  AOI211X1 U8352 ( .A0(n5073), .A1(n5478), .B0(n7298), .C0(n3357), .Y(n7291)
         );
  CLKINVX1 U8353 ( .A(n4881), .Y(n7302) );
  CLKINVX1 U8354 ( .A(n7305), .Y(n7301) );
  CLKINVX1 U8355 ( .A(n7300), .Y(n7297) );
  NAND2X1 U8356 ( .A(n7309), .B(n7204), .Y(n7305) );
  OAI21XL U8357 ( .A0(n7312), .A1(n5484), .B0(n7313), .Y(n8546) );
  MXI2X1 U8358 ( .A(\ImageBuffer[55][0] ), .B(n5039), .S0(n4882), .Y(n7313) );
  AOI211X1 U8359 ( .A0(n5073), .A1(n5487), .B0(n7320), .C0(n3357), .Y(n7312)
         );
  CLKINVX1 U8360 ( .A(n7322), .Y(n7319) );
  NAND2X1 U8361 ( .A(n7331), .B(n7203), .Y(n7327) );
  OAI21XL U8362 ( .A0(n7332), .A1(n5493), .B0(n7333), .Y(n8547) );
  AOI211X1 U8363 ( .A0(n7317), .A1(n7210), .B0(n7335), .C0(n7336), .Y(n7334)
         );
  AOI211X1 U8364 ( .A0(n5073), .A1(n5496), .B0(n7337), .C0(n3357), .Y(n7332)
         );
  OAI32X1 U8365 ( .A0(n7339), .A1(n7192), .A2(n7335), .B0(n5065), .B1(n7323), 
        .Y(n7338) );
  CLKINVX1 U8366 ( .A(n7339), .Y(n7336) );
  NAND2X1 U8367 ( .A(n7331), .B(n3396), .Y(n7342) );
  OAI21XL U8368 ( .A0(n7343), .A1(n5502), .B0(n7344), .Y(n8548) );
  MXI2X1 U8369 ( .A(\ImageBuffer[53][0] ), .B(n5039), .S0(n4884), .Y(n7344) );
  AOI211X1 U8370 ( .A0(n5073), .A1(n5505), .B0(n7348), .C0(n3358), .Y(n7343)
         );
  CLKINVX1 U8371 ( .A(n7350), .Y(n7347) );
  NAND2X1 U8372 ( .A(n7331), .B(n7235), .Y(n7353) );
  OAI21XL U8373 ( .A0(n7355), .A1(n5511), .B0(n7356), .Y(n8549) );
  OAI222XL U8374 ( .A0(n5516), .A1(n5045), .B0(n5517), .B1(n5048), .C0(n5518), 
        .C1(n5050), .Y(n7360) );
  OAI32X1 U8375 ( .A0(n7362), .A1(n7192), .A2(n7358), .B0(n5067), .B1(n7323), 
        .Y(n7361) );
  CLKINVX1 U8376 ( .A(n7362), .Y(n7359) );
  OAI21XL U8377 ( .A0(n7366), .A1(n5520), .B0(n7367), .Y(n8550) );
  AOI211X1 U8378 ( .A0(n7317), .A1(n7255), .B0(n7369), .C0(n7370), .Y(n7368)
         );
  AOI211X1 U8379 ( .A0(n5073), .A1(n5523), .B0(n7371), .C0(n3358), .Y(n7366)
         );
  OAI222XL U8380 ( .A0(n5525), .A1(n5045), .B0(n5526), .B1(n5048), .C0(n5527), 
        .C1(n5050), .Y(n7371) );
  OAI32X1 U8381 ( .A0(n7373), .A1(n7192), .A2(n7369), .B0(n3560), .B1(n7323), 
        .Y(n7372) );
  CLKINVX1 U8382 ( .A(n7373), .Y(n7370) );
  NAND2X1 U8383 ( .A(n7331), .B(n3397), .Y(n7376) );
  OAI21XL U8384 ( .A0(n7377), .A1(n5529), .B0(n7378), .Y(n8551) );
  MXI2X1 U8385 ( .A(\ImageBuffer[50][0] ), .B(n5039), .S0(n4887), .Y(n7378) );
  AOI211X1 U8386 ( .A0(n5073), .A1(n5532), .B0(n7382), .C0(n7187), .Y(n7377)
         );
  CLKINVX1 U8387 ( .A(n7384), .Y(n7381) );
  NAND2X1 U8388 ( .A(n7331), .B(n7277), .Y(n7387) );
  OAI21XL U8389 ( .A0(n7389), .A1(n5538), .B0(n7390), .Y(n8552) );
  OAI222XL U8390 ( .A0(n5543), .A1(n5045), .B0(n5544), .B1(n5048), .C0(n5545), 
        .C1(n5050), .Y(n7394) );
  OAI32X1 U8391 ( .A0(n7396), .A1(n7192), .A2(n7392), .B0(n5070), .B1(n7323), 
        .Y(n7395) );
  CLKINVX1 U8392 ( .A(n7396), .Y(n7393) );
  OAI21XL U8393 ( .A0(n7400), .A1(n5547), .B0(n7401), .Y(n8553) );
  AOI211X1 U8394 ( .A0(n7317), .A1(n7295), .B0(n7403), .C0(n7404), .Y(n7402)
         );
  AOI211X1 U8395 ( .A0(n5073), .A1(n5550), .B0(n7406), .C0(n7187), .Y(n7400)
         );
  OAI222XL U8396 ( .A0(n5552), .A1(n5045), .B0(n5553), .B1(n5048), .C0(n5554), 
        .C1(n5050), .Y(n7406) );
  OAI33X1 U8397 ( .A0(n7408), .A1(n7192), .A2(n7403), .B0(n7323), .B1(n7409), 
        .B2(n5071), .Y(n7407) );
  CLKINVX1 U8398 ( .A(n7412), .Y(n7409) );
  CLKINVX1 U8399 ( .A(n4890), .Y(n7410) );
  CLKINVX1 U8400 ( .A(n7408), .Y(n7404) );
  NAND2X1 U8401 ( .A(n7331), .B(n7309), .Y(n7412) );
  OAI21XL U8402 ( .A0(n7414), .A1(n5556), .B0(n7415), .Y(n8554) );
  MXI2X1 U8403 ( .A(\ImageBuffer[47][0] ), .B(n5038), .S0(n4891), .Y(n7415) );
  AOI211X1 U8404 ( .A0(n5073), .A1(n5559), .B0(n7421), .C0(n3358), .Y(n7414)
         );
  CLKINVX1 U8405 ( .A(n7423), .Y(n7420) );
  NAND2X1 U8406 ( .A(n7431), .B(n7203), .Y(n7427) );
  OAI21XL U8407 ( .A0(n7432), .A1(n5565), .B0(n7433), .Y(n8555) );
  AOI211X1 U8408 ( .A0(n7418), .A1(n7210), .B0(n7435), .C0(n7436), .Y(n7434)
         );
  AOI211X1 U8409 ( .A0(n5073), .A1(n5568), .B0(n7437), .C0(n3357), .Y(n7432)
         );
  OAI222XL U8410 ( .A0(n5570), .A1(n5045), .B0(n5571), .B1(n5047), .C0(n5572), 
        .C1(n5049), .Y(n7437) );
  OAI32X1 U8411 ( .A0(n7439), .A1(n7192), .A2(n7435), .B0(n3547), .B1(n3367), 
        .Y(n7438) );
  CLKINVX1 U8412 ( .A(n7439), .Y(n7436) );
  OAI21XL U8413 ( .A0(n7443), .A1(n5574), .B0(n7444), .Y(n8556) );
  MXI2X1 U8414 ( .A(\ImageBuffer[45][0] ), .B(n5038), .S0(n4893), .Y(n7444) );
  AOI211X1 U8415 ( .A0(n7418), .A1(n7224), .B0(n7446), .C0(n7447), .Y(n7445)
         );
  AOI211X1 U8416 ( .A0(n5073), .A1(n5577), .B0(n7448), .C0(n7187), .Y(n7443)
         );
  CLKINVX1 U8417 ( .A(n7450), .Y(n7447) );
  NAND2X1 U8418 ( .A(n7431), .B(n7235), .Y(n7453) );
  OAI21XL U8419 ( .A0(n7455), .A1(n5583), .B0(n7456), .Y(n8557) );
  OAI222XL U8420 ( .A0(n5588), .A1(n5045), .B0(n5589), .B1(n5047), .C0(n5590), 
        .C1(n5050), .Y(n7460) );
  OAI32X1 U8421 ( .A0(n7462), .A1(n7192), .A2(n7458), .B0(n3549), .B1(n3367), 
        .Y(n7461) );
  CLKINVX1 U8422 ( .A(n7462), .Y(n7459) );
  NAND2X1 U8423 ( .A(n7431), .B(n7250), .Y(n7465) );
  OAI21XL U8424 ( .A0(n7466), .A1(n5592), .B0(n7467), .Y(n8558) );
  OAI222XL U8425 ( .A0(n5597), .A1(n5045), .B0(n5598), .B1(n5047), .C0(n5599), 
        .C1(n5050), .Y(n7471) );
  OAI32X1 U8426 ( .A0(n7473), .A1(n7192), .A2(n7469), .B0(n5068), .B1(n3367), 
        .Y(n7472) );
  CLKINVX1 U8427 ( .A(n7473), .Y(n7470) );
  NAND2X1 U8428 ( .A(n7431), .B(n3397), .Y(n7476) );
  OAI21XL U8429 ( .A0(n7477), .A1(n5601), .B0(n7478), .Y(n8559) );
  MXI2X1 U8430 ( .A(\ImageBuffer[42][0] ), .B(n5038), .S0(n4896), .Y(n7478) );
  AOI211X1 U8431 ( .A0(n5073), .A1(n5604), .B0(n7482), .C0(n3357), .Y(n7477)
         );
  CLKINVX1 U8432 ( .A(n7484), .Y(n7481) );
  NAND2X1 U8433 ( .A(n7431), .B(n7277), .Y(n7487) );
  OAI21XL U8434 ( .A0(n7489), .A1(n5610), .B0(n7490), .Y(n8560) );
  OAI32X1 U8435 ( .A0(n7496), .A1(n7192), .A2(n7492), .B0(n5070), .B1(n3367), 
        .Y(n7495) );
  CLKINVX1 U8436 ( .A(n7496), .Y(n7493) );
  OAI21XL U8437 ( .A0(n7500), .A1(n5619), .B0(n7501), .Y(n8561) );
  OAI222XL U8438 ( .A0(n5624), .A1(n5045), .B0(n5625), .B1(n5047), .C0(n5626), 
        .C1(n5050), .Y(n7507) );
  OAI33X1 U8439 ( .A0(n7509), .A1(n7192), .A2(n7503), .B0(n3367), .B1(n7510), 
        .B2(n5071), .Y(n7508) );
  CLKINVX1 U8440 ( .A(n7513), .Y(n7510) );
  CLKINVX1 U8441 ( .A(n4899), .Y(n7511) );
  CLKINVX1 U8442 ( .A(n7509), .Y(n7504) );
  NAND2X1 U8443 ( .A(n7431), .B(n7309), .Y(n7513) );
  OAI21XL U8444 ( .A0(n7516), .A1(n5628), .B0(n7517), .Y(n8562) );
  MXI2X1 U8445 ( .A(\ImageBuffer[39][0] ), .B(n5038), .S0(n4900), .Y(n7517) );
  AOI211X1 U8446 ( .A0(n5073), .A1(n5631), .B0(n7523), .C0(n7187), .Y(n7516)
         );
  CLKINVX1 U8447 ( .A(n7525), .Y(n7522) );
  NAND2X1 U8448 ( .A(n7534), .B(n7203), .Y(n7530) );
  OAI21XL U8449 ( .A0(n7535), .A1(n5637), .B0(n7536), .Y(n8563) );
  AOI211X1 U8450 ( .A0(n7520), .A1(n7210), .B0(n7538), .C0(n7539), .Y(n7537)
         );
  OAI222XL U8451 ( .A0(n5642), .A1(n5045), .B0(n5643), .B1(n5047), .C0(n5644), 
        .C1(n5050), .Y(n7540) );
  OAI32X1 U8452 ( .A0(n7542), .A1(n7192), .A2(n7538), .B0(n5065), .B1(n7526), 
        .Y(n7541) );
  CLKINVX1 U8453 ( .A(n7542), .Y(n7539) );
  NAND2X1 U8454 ( .A(n7534), .B(n3396), .Y(n7545) );
  OAI21XL U8455 ( .A0(n7546), .A1(n5646), .B0(n7547), .Y(n8564) );
  MXI2X1 U8456 ( .A(\ImageBuffer[37][0] ), .B(n5038), .S0(n4902), .Y(n7547) );
  AOI211X1 U8457 ( .A0(n5073), .A1(n5649), .B0(n7551), .C0(n3358), .Y(n7546)
         );
  CLKINVX1 U8458 ( .A(n7553), .Y(n7550) );
  NAND2X1 U8459 ( .A(n7534), .B(n7235), .Y(n7556) );
  OAI21XL U8460 ( .A0(n7558), .A1(n5655), .B0(n7559), .Y(n8565) );
  OAI222XL U8461 ( .A0(n5660), .A1(n5045), .B0(n5661), .B1(n5047), .C0(n5662), 
        .C1(n5050), .Y(n7563) );
  OAI32X1 U8462 ( .A0(n7565), .A1(n7192), .A2(n7561), .B0(n5067), .B1(n7526), 
        .Y(n7564) );
  CLKINVX1 U8463 ( .A(n7565), .Y(n7562) );
  NAND2X1 U8464 ( .A(n7534), .B(n7250), .Y(n7568) );
  OAI21XL U8465 ( .A0(n7569), .A1(n5664), .B0(n7570), .Y(n8566) );
  AOI211X1 U8466 ( .A0(n7520), .A1(n7255), .B0(n7572), .C0(n7573), .Y(n7571)
         );
  OAI222XL U8467 ( .A0(n5669), .A1(n5045), .B0(n5670), .B1(n5048), .C0(n5671), 
        .C1(n5050), .Y(n7574) );
  OAI32X1 U8468 ( .A0(n7576), .A1(n7192), .A2(n7572), .B0(n5068), .B1(n7526), 
        .Y(n7575) );
  CLKINVX1 U8469 ( .A(n7576), .Y(n7573) );
  OAI21XL U8470 ( .A0(n7580), .A1(n5673), .B0(n7581), .Y(n8567) );
  MXI2X1 U8471 ( .A(\ImageBuffer[34][0] ), .B(n5040), .S0(n4905), .Y(n7581) );
  AOI211X1 U8472 ( .A0(n5073), .A1(n5676), .B0(n7585), .C0(n7187), .Y(n7580)
         );
  CLKINVX1 U8473 ( .A(n7587), .Y(n7584) );
  NAND2X1 U8474 ( .A(n7534), .B(n7277), .Y(n7590) );
  OAI21XL U8475 ( .A0(n7592), .A1(n5682), .B0(n7593), .Y(n8568) );
  AOI211X1 U8476 ( .A0(n7520), .A1(n7282), .B0(n7595), .C0(n7596), .Y(n7594)
         );
  OAI222XL U8477 ( .A0(n5687), .A1(n5045), .B0(n5688), .B1(n5047), .C0(n5689), 
        .C1(n5050), .Y(n7597) );
  CLKINVX1 U8478 ( .A(n7599), .Y(n7596) );
  MXI2X1 U8479 ( .A(\ImageBuffer[32][0] ), .B(n5038), .S0(n4907), .Y(n7604) );
  OAI222XL U8480 ( .A0(n5696), .A1(n5046), .B0(n5697), .B1(n5047), .C0(n5698), 
        .C1(n5050), .Y(n7608) );
  CLKINVX1 U8481 ( .A(n7614), .Y(n7611) );
  CLKINVX1 U8482 ( .A(n4908), .Y(n7612) );
  CLKINVX1 U8483 ( .A(n7610), .Y(n7607) );
  NAND2X1 U8484 ( .A(n7534), .B(n7309), .Y(n7614) );
  OAI21XL U8485 ( .A0(n7616), .A1(n5700), .B0(n7617), .Y(n8570) );
  MXI2X1 U8486 ( .A(\ImageBuffer[31][0] ), .B(n5038), .S0(n4909), .Y(n7617) );
  AOI211X1 U8487 ( .A0(n5073), .A1(n5703), .B0(n7623), .C0(n7187), .Y(n7616)
         );
  NAND2X1 U8488 ( .A(n7632), .B(n7200), .Y(n7625) );
  NAND2X1 U8489 ( .A(n7634), .B(n7203), .Y(n7630) );
  AOI211X1 U8490 ( .A0(n7620), .A1(n7210), .B0(n7638), .C0(n7639), .Y(n7637)
         );
  OAI32X1 U8491 ( .A0(n7642), .A1(n7192), .A2(n7638), .B0(n5065), .B1(n4825), 
        .Y(n7641) );
  NAND2X1 U8492 ( .A(n7634), .B(n3396), .Y(n7645) );
  OAI21XL U8493 ( .A0(n7646), .A1(n5718), .B0(n7647), .Y(n8572) );
  MXI2X1 U8494 ( .A(\ImageBuffer[29][0] ), .B(n5039), .S0(n4911), .Y(n7647) );
  AOI211X1 U8495 ( .A0(n5073), .A1(n5721), .B0(n7651), .C0(n3357), .Y(n7646)
         );
  NAND2X1 U8496 ( .A(n7632), .B(n7234), .Y(n7653) );
  NAND2X1 U8497 ( .A(n7634), .B(n7235), .Y(n7656) );
  OAI21XL U8498 ( .A0(n7658), .A1(n5727), .B0(n7659), .Y(n8573) );
  AOI211X1 U8499 ( .A0(n7620), .A1(n7240), .B0(n7661), .C0(n7662), .Y(n7660)
         );
  OAI32X1 U8500 ( .A0(n7665), .A1(n7192), .A2(n7661), .B0(n3549), .B1(n4825), 
        .Y(n7664) );
  NAND2X1 U8501 ( .A(n7634), .B(n7250), .Y(n7668) );
  OAI222XL U8502 ( .A0(n5741), .A1(n5046), .B0(n5742), .B1(n5047), .C0(n5743), 
        .C1(n5050), .Y(n7674) );
  OAI21XL U8503 ( .A0(n7680), .A1(n5745), .B0(n7681), .Y(n8575) );
  MXI2X1 U8504 ( .A(\ImageBuffer[26][0] ), .B(n5040), .S0(n4914), .Y(n7681) );
  AOI211X1 U8505 ( .A0(n5072), .A1(n5748), .B0(n7685), .C0(n7187), .Y(n7680)
         );
  NAND2X1 U8506 ( .A(n7634), .B(n7277), .Y(n7690) );
  OAI21XL U8507 ( .A0(n7692), .A1(n5754), .B0(n7693), .Y(n8576) );
  OAI32X1 U8508 ( .A0(n7699), .A1(n7192), .A2(n7695), .B0(n3559), .B1(n4825), 
        .Y(n7698) );
  OAI21XL U8509 ( .A0(n7703), .A1(n5763), .B0(n7704), .Y(n8577) );
  OAI222XL U8510 ( .A0(n5768), .A1(n5045), .B0(n5769), .B1(n5047), .C0(n5770), 
        .C1(n5050), .Y(n7709) );
  OAI33X1 U8511 ( .A0(n7711), .A1(n7192), .A2(n7706), .B0(n4825), .B1(n7712), 
        .B2(n5071), .Y(n7710) );
  CLKINVX1 U8512 ( .A(n7715), .Y(n7712) );
  CLKINVX1 U8513 ( .A(n4917), .Y(n7713) );
  NAND2X1 U8514 ( .A(n7634), .B(n7309), .Y(n7715) );
  OAI21XL U8515 ( .A0(n7718), .A1(n5772), .B0(n7719), .Y(n8578) );
  MXI2X1 U8516 ( .A(\ImageBuffer[23][0] ), .B(n5040), .S0(n4918), .Y(n7719) );
  AOI211X1 U8517 ( .A0(n5072), .A1(n5775), .B0(n7725), .C0(n7187), .Y(n7718)
         );
  NAND2X1 U8518 ( .A(n7735), .B(n7203), .Y(n7731) );
  OAI21XL U8519 ( .A0(n7736), .A1(n5781), .B0(n7737), .Y(n8579) );
  MXI2X1 U8520 ( .A(\ImageBuffer[22][0] ), .B(n5040), .S0(n4919), .Y(n7737) );
  AOI211X1 U8521 ( .A0(n7722), .A1(n7210), .B0(n7739), .C0(n7740), .Y(n7738)
         );
  AOI211X1 U8522 ( .A0(n5072), .A1(n5784), .B0(n7741), .C0(n3357), .Y(n7736)
         );
  NAND2X1 U8523 ( .A(n7733), .B(n7219), .Y(n7743) );
  OAI21XL U8524 ( .A0(n7747), .A1(n5790), .B0(n7748), .Y(n8580) );
  MXI2X1 U8525 ( .A(\ImageBuffer[21][0] ), .B(n5040), .S0(n4920), .Y(n7748) );
  AOI211X1 U8526 ( .A0(n5072), .A1(n5793), .B0(n7752), .C0(n3358), .Y(n7747)
         );
  NAND2X1 U8527 ( .A(n7735), .B(n7235), .Y(n7757) );
  OAI21XL U8528 ( .A0(n7759), .A1(n5799), .B0(n7760), .Y(n8581) );
  MXI2X1 U8529 ( .A(\ImageBuffer[20][0] ), .B(n5040), .S0(n4921), .Y(n7760) );
  AOI211X1 U8530 ( .A0(n7722), .A1(n7240), .B0(n7762), .C0(n7763), .Y(n7761)
         );
  AOI211X1 U8531 ( .A0(n5072), .A1(n5802), .B0(n7764), .C0(n3358), .Y(n7759)
         );
  NAND2X1 U8532 ( .A(n7733), .B(n7249), .Y(n7766) );
  NAND2X1 U8533 ( .A(n7735), .B(n7250), .Y(n7769) );
  OAI21XL U8534 ( .A0(n7770), .A1(n5808), .B0(n7771), .Y(n8582) );
  MXI2X1 U8535 ( .A(\ImageBuffer[19][0] ), .B(n5040), .S0(n4922), .Y(n7771) );
  AOI211X1 U8536 ( .A0(n5072), .A1(n5811), .B0(n7775), .C0(n7187), .Y(n7770)
         );
  OAI222XL U8537 ( .A0(n5813), .A1(n5045), .B0(n5814), .B1(n5047), .C0(n5815), 
        .C1(n5050), .Y(n7775) );
  NAND2X1 U8538 ( .A(n7735), .B(n3397), .Y(n7780) );
  OAI21XL U8539 ( .A0(n7781), .A1(n5817), .B0(n7782), .Y(n8583) );
  MXI2X1 U8540 ( .A(\ImageBuffer[18][0] ), .B(n5040), .S0(n4923), .Y(n7782) );
  AOI211X1 U8541 ( .A0(n5072), .A1(n5820), .B0(n7786), .C0(n7187), .Y(n7781)
         );
  NAND2X1 U8542 ( .A(n7735), .B(n7277), .Y(n7791) );
  OAI21XL U8543 ( .A0(n7793), .A1(n5826), .B0(n7794), .Y(n8584) );
  MXI2X1 U8544 ( .A(\ImageBuffer[17][0] ), .B(n5039), .S0(n4924), .Y(n7794) );
  AOI211X1 U8545 ( .A0(n5072), .A1(n5829), .B0(n7798), .C0(n3357), .Y(n7793)
         );
  MXI2X1 U8546 ( .A(\ImageBuffer[16][0] ), .B(n5038), .S0(n4925), .Y(n7805) );
  OAI222XL U8547 ( .A0(n5840), .A1(n5045), .B0(n5841), .B1(n5047), .C0(n5842), 
        .C1(n7189), .Y(n7809) );
  CLKINVX1 U8548 ( .A(n7815), .Y(n7812) );
  CLKINVX1 U8549 ( .A(n4926), .Y(n7813) );
  CLKINVX1 U8550 ( .A(n7811), .Y(n7808) );
  NAND2X1 U8551 ( .A(n7735), .B(n7309), .Y(n7815) );
  NAND3X1 U8552 ( .A(n5127), .B(n7717), .C(N2497), .Y(n7734) );
  OAI21XL U8553 ( .A0(n7817), .A1(n5844), .B0(n7818), .Y(n8586) );
  MXI2X1 U8554 ( .A(\ImageBuffer[15][0] ), .B(n5040), .S0(n4927), .Y(n7818) );
  AOI211X1 U8555 ( .A0(n7821), .A1(n7182), .B0(n7822), .C0(n7823), .Y(n7820)
         );
  AOI211X1 U8556 ( .A0(n5072), .A1(n5847), .B0(n7824), .C0(n3358), .Y(n7817)
         );
  CLKINVX1 U8557 ( .A(n7830), .Y(n7827) );
  NAND2X1 U8558 ( .A(n7832), .B(n7200), .Y(n7826) );
  NAND2X1 U8559 ( .A(n7834), .B(n7203), .Y(n7830) );
  OAI21XL U8560 ( .A0(n7835), .A1(n5853), .B0(n7836), .Y(n8587) );
  MXI2X1 U8561 ( .A(\ImageBuffer[14][0] ), .B(n5038), .S0(n4928), .Y(n7836) );
  AOI211X1 U8562 ( .A0(n7821), .A1(n7210), .B0(n7838), .C0(n7839), .Y(n7837)
         );
  OAI32X1 U8563 ( .A0(n7838), .A1(n5058), .A2(n7839), .B0(n3352), .B1(n7845), 
        .Y(n7844) );
  OAI21XL U8564 ( .A0(n7846), .A1(n5862), .B0(n7847), .Y(n8588) );
  MXI2X1 U8565 ( .A(\ImageBuffer[13][0] ), .B(n5040), .S0(n4929), .Y(n7847) );
  AOI211X1 U8566 ( .A0(n5072), .A1(n5865), .B0(n7851), .C0(n7187), .Y(n7846)
         );
  CLKINVX1 U8567 ( .A(n7856), .Y(n7854) );
  NAND2X1 U8568 ( .A(n7832), .B(n7234), .Y(n7853) );
  NAND2X1 U8569 ( .A(n7834), .B(n7235), .Y(n7856) );
  OAI21XL U8570 ( .A0(n7858), .A1(n5871), .B0(n7859), .Y(n8589) );
  MXI2X1 U8571 ( .A(\ImageBuffer[12][0] ), .B(n5040), .S0(n4930), .Y(n7859) );
  OAI32X1 U8572 ( .A0(n7861), .A1(n5058), .A2(n7862), .B0(n3351), .B1(n7868), 
        .Y(n7867) );
  OAI21XL U8573 ( .A0(n7869), .A1(n5880), .B0(n7870), .Y(n8590) );
  AOI211X1 U8574 ( .A0(n5072), .A1(n5883), .B0(n7874), .C0(n3358), .Y(n7869)
         );
  OAI222XL U8575 ( .A0(n5885), .A1(n5046), .B0(n5886), .B1(n5048), .C0(n5887), 
        .C1(n5049), .Y(n7874) );
  OAI32X1 U8576 ( .A0(n7876), .A1(n7192), .A2(n7872), .B0(n5068), .B1(n3369), 
        .Y(n7875) );
  OAI21XL U8577 ( .A0(n7880), .A1(n5889), .B0(n7881), .Y(n8591) );
  MXI2X1 U8578 ( .A(\ImageBuffer[10][0] ), .B(n5040), .S0(n4932), .Y(n7881) );
  CLKINVX1 U8579 ( .A(n7890), .Y(n7888) );
  NAND2X1 U8580 ( .A(n7834), .B(n7277), .Y(n7890) );
  OAI21XL U8581 ( .A0(n7892), .A1(n5898), .B0(n7893), .Y(n8592) );
  AOI211X1 U8582 ( .A0(n5072), .A1(n5901), .B0(n7897), .C0(n3358), .Y(n7892)
         );
  OAI222XL U8583 ( .A0(n5903), .A1(n5046), .B0(n5904), .B1(n5048), .C0(n5905), 
        .C1(n5049), .Y(n7897) );
  OAI21XL U8584 ( .A0(n7903), .A1(n5907), .B0(n7904), .Y(n8593) );
  AOI211X1 U8585 ( .A0(n5072), .A1(n5910), .B0(n7908), .C0(n7187), .Y(n7903)
         );
  OAI222XL U8586 ( .A0(n5912), .A1(n5046), .B0(n5913), .B1(n5048), .C0(n5914), 
        .C1(n5049), .Y(n7908) );
  CLKINVX1 U8587 ( .A(n7914), .Y(n7911) );
  CLKINVX1 U8588 ( .A(n7833), .Y(n7912) );
  OAI32X1 U8589 ( .A0(n7906), .A1(n5058), .A2(n7907), .B0(n3351), .B1(n7914), 
        .Y(n7915) );
  NAND2X1 U8590 ( .A(n7834), .B(n7309), .Y(n7914) );
  OAI21XL U8591 ( .A0(n7916), .A1(n5916), .B0(n7917), .Y(n8594) );
  MXI2X1 U8592 ( .A(\ImageBuffer[7][0] ), .B(n5039), .S0(n4935), .Y(n7917) );
  AOI211X1 U8593 ( .A0(n7182), .A1(n3371), .B0(n7920), .C0(n7921), .Y(n7919)
         );
  NAND2X1 U8594 ( .A(n7923), .B(n7924), .Y(n7315) );
  CLKINVX1 U8595 ( .A(n7932), .Y(n7929) );
  NAND2X1 U8596 ( .A(n7934), .B(n7200), .Y(n7927) );
  NAND2X1 U8597 ( .A(n7936), .B(n7203), .Y(n7932) );
  OAI21XL U8598 ( .A0(n7937), .A1(n5925), .B0(n7938), .Y(n8595) );
  MXI2X1 U8599 ( .A(\ImageBuffer[6][0] ), .B(n5040), .S0(n4936), .Y(n7938) );
  AOI211X1 U8600 ( .A0(n5072), .A1(n5928), .B0(n7943), .C0(n3357), .Y(n7937)
         );
  OAI21XL U8601 ( .A0(n7949), .A1(n5934), .B0(n7950), .Y(n8596) );
  MXI2X1 U8602 ( .A(\ImageBuffer[5][0] ), .B(n7178), .S0(n4937), .Y(n7950) );
  AOI211X1 U8603 ( .A0(n5072), .A1(n5937), .B0(n7955), .C0(n3358), .Y(n7949)
         );
  CLKINVX1 U8604 ( .A(n7960), .Y(n7958) );
  NAND2X1 U8605 ( .A(n7936), .B(n7235), .Y(n7960) );
  OAI21XL U8606 ( .A0(n7962), .A1(n5943), .B0(n7963), .Y(n8597) );
  MXI2X1 U8607 ( .A(\ImageBuffer[4][0] ), .B(n7178), .S0(n4938), .Y(n7963) );
  NOR2X1 U8608 ( .A(n4945), .B(n7968), .Y(n7923) );
  AOI211X1 U8609 ( .A0(n5072), .A1(n5946), .B0(n7969), .C0(n7187), .Y(n7962)
         );
  OAI21XL U8610 ( .A0(n7975), .A1(n5952), .B0(n7976), .Y(n8598) );
  MXI2X1 U8611 ( .A(\ImageBuffer[3][0] ), .B(n5039), .S0(n4939), .Y(n7976) );
  AOI211X1 U8612 ( .A0(n5072), .A1(n5955), .B0(n7981), .C0(n3357), .Y(n7975)
         );
  NAND2X1 U8613 ( .A(n7934), .B(n3395), .Y(n7983) );
  NOR2X1 U8614 ( .A(n5117), .B(n3935), .Y(n7922) );
  OAI21XL U8615 ( .A0(n7987), .A1(n5961), .B0(n7988), .Y(n8599) );
  AOI211X1 U8616 ( .A0(n5072), .A1(n5964), .B0(n7992), .C0(n7187), .Y(n7987)
         );
  OAI222XL U8617 ( .A0(n5966), .A1(n5046), .B0(n5967), .B1(n5047), .C0(n5968), 
        .C1(n5049), .Y(n7992) );
  OAI33X1 U8618 ( .A0(n7994), .A1(n7192), .A2(n7990), .B0(n7928), .B1(n7995), 
        .B2(n5069), .Y(n7993) );
  OAI33X1 U8619 ( .A0(n7994), .A1(n5053), .A2(n7990), .B0(n7931), .B1(n7995), 
        .B2(n5069), .Y(n7996) );
  CLKINVX1 U8620 ( .A(n7997), .Y(n7995) );
  NAND2X1 U8621 ( .A(n7936), .B(n7277), .Y(n7997) );
  OAI21XL U8622 ( .A0(n7999), .A1(n5970), .B0(n8000), .Y(n8600) );
  MXI2X1 U8623 ( .A(\ImageBuffer[1][0] ), .B(n5038), .S0(n4941), .Y(n8000) );
  AOI211X1 U8624 ( .A0(n5072), .A1(n5973), .B0(n8004), .C0(n3358), .Y(n7999)
         );
  OAI21XL U8625 ( .A0(n8010), .A1(n5979), .B0(n8011), .Y(n8601) );
  MXI2X1 U8626 ( .A(\ImageBuffer[0][0] ), .B(n5040), .S0(n4942), .Y(n8011) );
  NOR2BX1 U8627 ( .AN(IROM_Q[0]), .B(n4945), .Y(n7178) );
  NAND3BX1 U8628 ( .AN(n4943), .B(n8014), .C(n8015), .Y(n8013) );
  AOI211X1 U8629 ( .A0(n3371), .A1(n7295), .B0(n8016), .C0(n8017), .Y(n8012)
         );
  NOR2X1 U8630 ( .A(n4945), .B(n8620), .Y(n7980) );
  CLKINVX1 U8631 ( .A(n8018), .Y(n7179) );
  AOI211X1 U8632 ( .A0(n5073), .A1(n5983), .B0(n8019), .C0(n7187), .Y(n8010)
         );
  NAND2X1 U8633 ( .A(n8021), .B(n5404), .Y(n8014) );
  CLKINVX1 U8634 ( .A(N2781), .Y(n7189) );
  CLKINVX1 U8635 ( .A(n8027), .Y(n8024) );
  CLKINVX1 U8636 ( .A(n7935), .Y(n8025) );
  CLKINVX1 U8637 ( .A(n8023), .Y(n8017) );
  NAND2X1 U8638 ( .A(n7936), .B(n7309), .Y(n8027) );
  NAND2X1 U8639 ( .A(n7967), .B(n5115), .Y(\sub_168_aco/B[0] ) );
  NOR2X1 U8640 ( .A(n5118), .B(n3751), .Y(n7967) );
  OAI2BB2XL U8641 ( .B0(n7942), .B1(n8035), .A0N(n7942), .A1N(n8036), .Y(n3338) );
  OAI2BB2XL U8642 ( .B0(n7708), .B1(n8035), .A0N(N2549), .A1N(n8036), .Y(n3337) );
  OAI2BB2XL U8643 ( .B0(n7954), .B1(n8035), .A0N(N2545), .A1N(n8036), .Y(n3336) );
  OAI2BB2XL U8644 ( .B0(n7968), .B1(n8035), .A0N(N2546), .A1N(n8036), .Y(n3335) );
  OAI2BB2XL U8645 ( .B0(n7405), .B1(n8035), .A0N(N2547), .A1N(n8036), .Y(n3334) );
  OAI2BB2XL U8646 ( .B0(n7506), .B1(n8035), .A0N(N2548), .A1N(n8036), .Y(n3333) );
  NOR2X1 U8647 ( .A(n7954), .B(n7942), .Y(n7924) );
  NAND2X1 U8648 ( .A(n8602), .B(n4945), .Y(n8035) );
  NAND4BX1 U8649 ( .AN(n8040), .B(N2522), .C(n5104), .D(N2521), .Y(n8039) );
  NAND3X1 U8650 ( .A(n5105), .B(n5106), .C(N2519), .Y(n8040) );
  OAI221XL U8651 ( .A0(n8041), .A1(n8042), .B0(n8043), .B1(n4298), .C0(n8602), 
        .Y(n3326) );
  AOI221XL U8652 ( .A0(n8044), .A1(n3935), .B0(n5118), .B1(n3475), .C0(n8045), 
        .Y(n8041) );
  AO22X1 U8653 ( .A0(N2630), .A1(n3476), .B0(n5118), .B1(n3477), .Y(n8045) );
  OAI221XL U8654 ( .A0(n8046), .A1(n8042), .B0(n8043), .B1(n5117), .C0(n8602), 
        .Y(n3325) );
  AOI221XL U8655 ( .A0(n8044), .A1(n3929), .B0(n3748), .B1(n3475), .C0(n8047), 
        .Y(n8046) );
  AO22X1 U8656 ( .A0(N2631), .A1(n3476), .B0(n4122), .B1(n3477), .Y(n8047) );
  OAI22XL U8657 ( .A0(n8043), .A1(n5115), .B0(n8048), .B1(n8042), .Y(n3324) );
  AOI221XL U8658 ( .A0(n8044), .A1(n3409), .B0(N2495), .B1(n3475), .C0(n8049), 
        .Y(n8048) );
  OAI221XL U8659 ( .A0(n8050), .A1(n8042), .B0(n8043), .B1(n5128), .C0(n8602), 
        .Y(n3323) );
  AOI221XL U8660 ( .A0(n8044), .A1(N2490), .B0(N2623), .B1(n3475), .C0(n8051), 
        .Y(n8050) );
  AO22X1 U8661 ( .A0(N2633), .A1(n3476), .B0(N2613), .B1(n3477), .Y(n8051) );
  OAI221XL U8662 ( .A0(n8052), .A1(n8042), .B0(n8043), .B1(n5126), .C0(n8602), 
        .Y(n3322) );
  AOI221XL U8663 ( .A0(n8044), .A1(N2491), .B0(N2624), .B1(n3475), .C0(n8053), 
        .Y(n8052) );
  OAI22XL U8664 ( .A0(n8043), .A1(n7505), .B0(n8054), .B1(n8042), .Y(n3321) );
  AOI221XL U8665 ( .A0(n8044), .A1(N2492), .B0(N2625), .B1(n3475), .C0(n8055), 
        .Y(n8054) );
  AO22X1 U8666 ( .A0(N2635), .A1(n3476), .B0(N2615), .B1(n3477), .Y(n8055) );
  NOR2X1 U8667 ( .A(n8056), .B(n7210), .Y(n8044) );
  OAI31XL U8668 ( .A0(n8042), .A1(n8057), .A2(n8056), .B0(n8059), .Y(n8058) );
  NAND3X1 U8669 ( .A(n3756), .B(n3939), .C(N2495), .Y(n8057) );
  NAND2X1 U8670 ( .A(n8059), .B(n8602), .Y(n8042) );
  NAND3X1 U8671 ( .A(n5404), .B(n5405), .C(cmd[2]), .Y(n8056) );
  NAND2X1 U8672 ( .A(\state_cs[0] ), .B(n5400), .Y(n8018) );
  NAND2X1 U8673 ( .A(n5400), .B(n4945), .Y(n8629) );
  NAND2X1 U8674 ( .A(n4947), .B(n5125), .Y(N2617) );
  CLKINVX1 U8675 ( .A(n4947), .Y(n7505) );
  AOI2BB2X1 U8676 ( .B0(n8079), .B1(N2495), .A0N(n3408), .A1N(n8080), .Y(n8083) );
  LCD_CTRL_DW01_add_5 add_2_root_add_0_root_add_207_3 ( .A({1'b0, 1'b0, n5099, 
        n5094, n5093, n5090, n5083, n5081, n5075, n5072}), .B({1'b0, 1'b0, 
        n4861, n4862, n4863, n4864, n4865, N2779, n4866, N2781}), .CI(1'b0), 
        .SUM({SYNOPSYS_UNCONNECTED__0, N2740, N2739, N2738, N2737, N2736, 
        N2735, N2734, N2733, N2732}) );
  LCD_CTRL_DW01_add_4 add_1_root_add_0_root_add_207_3 ( .A({1'b0, N2740, N2739, 
        N2738, N2737, N2736, N2735, N2734, N2733, N2732}), .B({1'b0, 1'b0, 
        N2766, N2767, N2768, N2769, N2770, N2771, N2772, N2773}), .CI(1'b0), 
        .SUM({n8613, n8612, n8611, n8610, n8609, n8608, n8607, n8606, n8605, 
        n8604}) );
  LCD_CTRL_DW01_add_3 add_0_root_add_0_root_add_207_3 ( .A({1'b0, 1'b0, n4867, 
        n4868, n4869, n4870, n4871, n4872, n4873, N2765}), .B({n8613, n8612, 
        n8611, n8610, n8609, n8608, n8607, n8606, n8605, n8604}), .CI(1'b0), 
        .SUM({sum, SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2}) );
  EDFFXL \IRAM_D_reg[7]  ( .D(N13064), .E(IRAM_valid), .CK(clk), .QN(n3406) );
  EDFFHQX1 \IRAM_D_reg[2]  ( .D(N13069), .E(IRAM_valid), .CK(clk), .Q(n8649)
         );
  INVXL U4426 ( .A(n8645), .Y(n8631) );
  INVX12 U4427 ( .A(n8631), .Y(IRAM_D[6]) );
  INVXL U4428 ( .A(n8646), .Y(n8633) );
  INVX12 U4429 ( .A(n8633), .Y(IRAM_D[5]) );
  INVXL U4430 ( .A(n8647), .Y(n8635) );
  INVX12 U4431 ( .A(n8635), .Y(IRAM_D[4]) );
  INVXL U4432 ( .A(n8648), .Y(n8637) );
  INVX12 U4433 ( .A(n8637), .Y(IRAM_D[3]) );
  INVXL U8682 ( .A(n8650), .Y(n8639) );
  INVX12 U8683 ( .A(n8639), .Y(IRAM_D[1]) );
  INVXL U8684 ( .A(n8651), .Y(n8641) );
  INVX12 U8685 ( .A(n8641), .Y(IRAM_D[0]) );
  INVXL U8686 ( .A(n8649), .Y(n8643) );
  INVX12 U8687 ( .A(n8643), .Y(IRAM_D[2]) );
endmodule

